module top ();
    lib lib_i ();
endmodule
