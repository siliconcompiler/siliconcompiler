// Name: Black Parrot Back-end (BE) Only
//
// Description: Back-end of a 64-bit RISC-V Core with Cache Coherence Directory.
//
// Top Module: bp_be_top
//
// GitHub: https://github.com/black-parrot/pre-alpha-release
//    commit: ceb22c57f269726a5fd99b722521cf7df9d3907c
//

module bsg_dff_reset_en_64_80000124
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69;
  reg [63:0] data_o;
  assign N3 = (N0)? 1'b1 : 
              (N69)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = reset_i;
  assign { N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                        (N69)? data_i : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N68 = ~reset_i;
  assign N69 = en_i & N68;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[63:0] } <= { N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4 };
    end 
  end


endmodule



module bsg_mux_width_p64_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [0:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1;
  assign data_o[63] = (N1)? data_i[63] : 
                      (N0)? data_i[127] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[62] = (N1)? data_i[62] : 
                      (N0)? data_i[126] : 1'b0;
  assign data_o[61] = (N1)? data_i[61] : 
                      (N0)? data_i[125] : 1'b0;
  assign data_o[60] = (N1)? data_i[60] : 
                      (N0)? data_i[124] : 1'b0;
  assign data_o[59] = (N1)? data_i[59] : 
                      (N0)? data_i[123] : 1'b0;
  assign data_o[58] = (N1)? data_i[58] : 
                      (N0)? data_i[122] : 1'b0;
  assign data_o[57] = (N1)? data_i[57] : 
                      (N0)? data_i[121] : 1'b0;
  assign data_o[56] = (N1)? data_i[56] : 
                      (N0)? data_i[120] : 1'b0;
  assign data_o[55] = (N1)? data_i[55] : 
                      (N0)? data_i[119] : 1'b0;
  assign data_o[54] = (N1)? data_i[54] : 
                      (N0)? data_i[118] : 1'b0;
  assign data_o[53] = (N1)? data_i[53] : 
                      (N0)? data_i[117] : 1'b0;
  assign data_o[52] = (N1)? data_i[52] : 
                      (N0)? data_i[116] : 1'b0;
  assign data_o[51] = (N1)? data_i[51] : 
                      (N0)? data_i[115] : 1'b0;
  assign data_o[50] = (N1)? data_i[50] : 
                      (N0)? data_i[114] : 1'b0;
  assign data_o[49] = (N1)? data_i[49] : 
                      (N0)? data_i[113] : 1'b0;
  assign data_o[48] = (N1)? data_i[48] : 
                      (N0)? data_i[112] : 1'b0;
  assign data_o[47] = (N1)? data_i[47] : 
                      (N0)? data_i[111] : 1'b0;
  assign data_o[46] = (N1)? data_i[46] : 
                      (N0)? data_i[110] : 1'b0;
  assign data_o[45] = (N1)? data_i[45] : 
                      (N0)? data_i[109] : 1'b0;
  assign data_o[44] = (N1)? data_i[44] : 
                      (N0)? data_i[108] : 1'b0;
  assign data_o[43] = (N1)? data_i[43] : 
                      (N0)? data_i[107] : 1'b0;
  assign data_o[42] = (N1)? data_i[42] : 
                      (N0)? data_i[106] : 1'b0;
  assign data_o[41] = (N1)? data_i[41] : 
                      (N0)? data_i[105] : 1'b0;
  assign data_o[40] = (N1)? data_i[40] : 
                      (N0)? data_i[104] : 1'b0;
  assign data_o[39] = (N1)? data_i[39] : 
                      (N0)? data_i[103] : 1'b0;
  assign data_o[38] = (N1)? data_i[38] : 
                      (N0)? data_i[102] : 1'b0;
  assign data_o[37] = (N1)? data_i[37] : 
                      (N0)? data_i[101] : 1'b0;
  assign data_o[36] = (N1)? data_i[36] : 
                      (N0)? data_i[100] : 1'b0;
  assign data_o[35] = (N1)? data_i[35] : 
                      (N0)? data_i[99] : 1'b0;
  assign data_o[34] = (N1)? data_i[34] : 
                      (N0)? data_i[98] : 1'b0;
  assign data_o[33] = (N1)? data_i[33] : 
                      (N0)? data_i[97] : 1'b0;
  assign data_o[32] = (N1)? data_i[32] : 
                      (N0)? data_i[96] : 1'b0;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[95] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[94] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[93] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[92] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[91] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[90] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[89] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[88] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[87] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[86] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[85] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[84] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[83] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[82] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[81] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[80] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[79] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[78] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[77] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[76] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[75] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[74] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[73] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[72] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[71] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[70] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[69] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[68] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[67] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[66] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[65] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[64] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_dff_en_width_p36
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [35:0] data_i;
  output [35:0] data_o;
  input clk_i;
  input en_i;
  reg [35:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[35:0] } <= { data_i[35:0] };
    end 
  end


endmodule



module bsg_dff_reset_en_width_p1
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6;
  reg [0:0] data_o;
  assign N3 = (N0)? 1'b1 : 
              (N6)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = reset_i;
  assign N4 = (N0)? 1'b0 : 
              (N6)? data_i[0] : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N5 = ~reset_i;
  assign N6 = en_i & N5;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[0:0] } <= { N4 };
    end 
  end


endmodule



module bp_be_director_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
(
  clk_i,
  reset_i,
  calc_status_i,
  expected_npc_o,
  fe_cmd_o,
  fe_cmd_v_o,
  fe_cmd_ready_i,
  chk_flush_fe_o,
  chk_dequeue_fe_o,
  chk_roll_fe_o
);

  input [301:0] calc_status_i;
  output [63:0] expected_npc_o;
  output [108:0] fe_cmd_o;
  input clk_i;
  input reset_i;
  input fe_cmd_ready_i;
  output fe_cmd_v_o;
  output chk_flush_fe_o;
  output chk_dequeue_fe_o;
  output chk_roll_fe_o;
  wire [63:0] expected_npc_o,npc_n,npc_r,ret_mux_o,miss_mux_o,br_mux_o,npc_plus4;
  wire [108:0] fe_cmd_o;
  wire fe_cmd_v_o,chk_flush_fe_o,chk_dequeue_fe_o,chk_roll_fe_o,N0,N1,N2,N3,N4,N5,
  npc_w_v,btaken_v,npc_mismatch_v,redirect_pending,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,net16566,net16567,net16568,net16569,net16570,net16571,
  net16572,net16573,net16574,net16575,net16576,net16577,net16578,net16579,net16580,
  net16581,net16582,net16583,net16584,net16585,net16586,net16587,net16588,net16589,
  net16590,net16591,net16592,net16593,net16594,net16595,net16596,net16597,net16598,
  net16599,net16600,net16601,net16602,net16603,net16604,net16605,net16606,net16607,
  net16608,net16609,net16610,net16611,net16612,net16613,net16614,net16615,net16616,
  net16617,net16618,net16619,net16620,net16621,net16622,net16623,net16624,
  net16625,net16626,net16627,net16628,net16629,net16630,net16631,net16632,net16633,
  net16634,net16635,net16636,net16637,net16638,net16639,net16640,net16641,net16642,
  net16643,net16644,net16645,net16646,net16647,net16648,net16649,net16650,net16651,
  net16652,net16653,net16654,net16655,net16656,net16657,net16658,net16659,net16660,
  net16661,net16662,net16663,net16664,net16665,net16666,net16667,net16668,net16669,
  net16670,net16671,net16672,net16673,net16674,net16675,net16676,net16677,net16678,
  net16679,net16680,net16681,net16682,net16683,net16684,net16685,net16686,net16687,
  net16688,net16689,net16690,net16691,net16692,net16693;
  wire [35:0] branch_metadata_fwd_r;
  assign fe_cmd_o[107] = 1'b0;
  assign chk_roll_fe_o = calc_status_i[3];

  bsg_dff_reset_en_64_80000124
  npc
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(npc_w_v),
    .data_i(npc_n),
    .data_o(npc_r)
  );


  bsg_mux_width_p64_els_p2
  exception_mux
  (
    .data_i({ ret_mux_o, miss_mux_o }),
    .sel_i(calc_status_i[2]),
    .data_o(npc_n)
  );


  bsg_mux_width_p64_els_p2
  miss_mux
  (
    .data_i({ calc_status_i[67:4], br_mux_o }),
    .sel_i(calc_status_i[3]),
    .data_o(miss_mux_o)
  );


  bsg_mux_width_p64_els_p2
  br_mux
  (
    .data_i({ calc_status_i[221:158], npc_plus4 }),
    .sel_i(btaken_v),
    .data_o(br_mux_o)
  );


  bsg_mux_width_p64_els_p2
  ret_mux
  (
    .data_i({ net16566, net16567, net16568, net16569, net16570, net16571, net16572, net16573, net16574, net16575, net16576, net16577, net16578, net16579, net16580, net16581, net16582, net16583, net16584, net16585, net16586, net16587, net16588, net16589, net16590, net16591, net16592, net16593, net16594, net16595, net16596, net16597, net16598, net16599, net16600, net16601, net16602, net16603, net16604, net16605, net16606, net16607, net16608, net16609, net16610, net16611, net16612, net16613, net16614, net16615, net16616, net16617, net16618, net16619, net16620, net16621, net16622, net16623, net16624, net16625, net16626, net16627, net16628, net16629, net16630, net16631, net16632, net16633, net16634, net16635, net16636, net16637, net16638, net16639, net16640, net16641, net16642, net16643, net16644, net16645, net16646, net16647, net16648, net16649, net16650, net16651, net16652, net16653, net16654, net16655, net16656, net16657, net16658, net16659, net16660, net16661, net16662, net16663, net16664, net16665, net16666, net16667, net16668, net16669, net16670, net16671, net16672, net16673, net16674, net16675, net16676, net16677, net16678, net16679, net16680, net16681, net16682, net16683, net16684, net16685, net16686, net16687, net16688, net16689, net16690, net16691, net16692, net16693 }),
    .sel_i(calc_status_i[1]),
    .data_o(ret_mux_o)
  );


  bsg_dff_en_width_p36
  branch_metadata_fwd_reg
  (
    .clk_i(clk_i),
    .data_i(calc_status_i[157:122]),
    .en_i(calc_status_i[119]),
    .data_o(branch_metadata_fwd_r)
  );

  assign npc_mismatch_v = expected_npc_o != calc_status_i[300:237];

  bsg_dff_reset_en_width_p1
  redirect_pending_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(calc_status_i[301]),
    .data_i(npc_mismatch_v),
    .data_o(redirect_pending)
  );

  assign N90 = ~fe_cmd_o[106];
  assign N91 = N90 | fe_cmd_o[108];
  assign N92 = ~N91;
  assign npc_plus4 = npc_r + { 1'b1, 1'b0, 1'b0 };
  assign expected_npc_o = (N0)? npc_n : 
                          (N1)? npc_r : 1'b0;
  assign N0 = N7;
  assign N1 = N6;
  assign { N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12 } = (N2)? calc_status_i[157:122] : 
                                                                                                                                                                                                  (N51)? branch_metadata_fwd_r : 1'b0;
  assign N2 = N50;
  assign N48 = ~calc_status_i[121];
  assign { N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52 } = (N2)? calc_status_i[157:122] : 
                                                                                                                                                                                                  (N51)? branch_metadata_fwd_r : 1'b0;
  assign { fe_cmd_o[108:108], fe_cmd_o[105:0] } = (N3)? { 1'b0, expected_npc_o, 1'b1, 1'b0, 1'b0, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N48, 1'b0, 1'b0 } : 
                                                  (N4)? { 1'b1, calc_status_i[300:237], N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N3 = N8;
  assign N4 = N9;
  assign fe_cmd_o[106] = (N3)? 1'b1 : 
                         (N89)? 1'b0 : 
                         (N5)? 1'b0 : 1'b0;
  assign N5 = 1'b0;
  assign fe_cmd_v_o = (N3)? N49 : 
                      (N4)? N88 : 
                      (N11)? 1'b0 : 1'b0;
  assign npc_w_v = calc_status_i[119] | calc_status_i[3];
  assign btaken_v = calc_status_i[222] & calc_status_i[120];
  assign N6 = ~npc_w_v;
  assign N7 = npc_w_v;
  assign chk_dequeue_fe_o = N93 & calc_status_i[0];
  assign N93 = ~calc_status_i[3];
  assign chk_flush_fe_o = fe_cmd_v_o & N92;
  assign N8 = calc_status_i[301] & npc_mismatch_v;
  assign N9 = N95 & calc_status_i[121];
  assign N95 = calc_status_i[301] & N94;
  assign N94 = ~npc_mismatch_v;
  assign N10 = N9 | N8;
  assign N11 = ~N10;
  assign N49 = N97 & N98;
  assign N97 = fe_cmd_ready_i & N96;
  assign N96 = ~calc_status_i[3];
  assign N98 = ~redirect_pending;
  assign N50 = calc_status_i[119];
  assign N51 = ~N50;
  assign N88 = N100 & N98;
  assign N100 = fe_cmd_ready_i & N99;
  assign N99 = ~calc_status_i[3];
  assign N89 = ~N8;

endmodule



module bp_be_detector_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
(
  clk_i,
  reset_i,
  calc_status_i,
  expected_npc_i,
  mmu_cmd_ready_i,
  chk_dispatch_v_o,
  chk_roll_o,
  chk_poison_isd_o,
  chk_poison_ex_o
);

  input [301:0] calc_status_i;
  input [63:0] expected_npc_i;
  input clk_i;
  input reset_i;
  input mmu_cmd_ready_i;
  output chk_dispatch_v_o;
  output chk_roll_o;
  output chk_poison_isd_o;
  output chk_poison_ex_o;
  wire chk_dispatch_v_o,chk_roll_o,chk_poison_isd_o,chk_poison_ex_o,N0,N1,N2,N3,N4,N5,
  data_haz_v,struct_haz_v,N6,mispredict_v,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,
  N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,
  N38,N39,N40,N41,N42,N43,N44;
  wire [2:0] rs1_match_vector,rs2_match_vector,frs1_data_haz_v,frs2_data_haz_v;
  wire [1:0] irs1_data_haz_v,irs2_data_haz_v;
  assign chk_roll_o = calc_status_i[3];
  assign N0 = calc_status_i[234:230] == calc_status_i[73:69];
  assign N1 = calc_status_i[227:223] == calc_status_i[73:69];
  assign N2 = calc_status_i[234:230] == calc_status_i[83:79];
  assign N3 = calc_status_i[227:223] == calc_status_i[83:79];
  assign N4 = calc_status_i[234:230] == calc_status_i[93:89];
  assign N5 = calc_status_i[227:223] == calc_status_i[93:89];
  assign N6 = calc_status_i[300:237] != expected_npc_i;
  assign N7 = calc_status_i[233] | calc_status_i[234];
  assign N8 = calc_status_i[232] | N7;
  assign N9 = calc_status_i[231] | N8;
  assign N10 = calc_status_i[230] | N9;
  assign N11 = calc_status_i[226] | calc_status_i[227];
  assign N12 = calc_status_i[225] | N11;
  assign N13 = calc_status_i[224] | N12;
  assign N14 = calc_status_i[223] | N13;
  assign rs1_match_vector[0] = N10 & N0;
  assign rs2_match_vector[0] = N14 & N1;
  assign rs1_match_vector[1] = N10 & N2;
  assign rs2_match_vector[1] = N14 & N3;
  assign rs1_match_vector[2] = N10 & N4;
  assign rs2_match_vector[2] = N14 & N5;
  assign irs1_data_haz_v[0] = N15 & N16;
  assign N15 = calc_status_i[236] & rs1_match_vector[0];
  assign N16 = calc_status_i[77] | calc_status_i[76];
  assign irs2_data_haz_v[0] = N17 & N18;
  assign N17 = calc_status_i[229] & rs2_match_vector[0];
  assign N18 = calc_status_i[77] | calc_status_i[76];
  assign frs1_data_haz_v[0] = N19 & N20;
  assign N19 = calc_status_i[235] & rs1_match_vector[0];
  assign N20 = calc_status_i[75] | calc_status_i[74];
  assign frs2_data_haz_v[0] = N21 & N22;
  assign N21 = calc_status_i[228] & rs2_match_vector[0];
  assign N22 = calc_status_i[75] | calc_status_i[74];
  assign irs1_data_haz_v[1] = N23 & calc_status_i[86];
  assign N23 = calc_status_i[236] & rs1_match_vector[1];
  assign irs2_data_haz_v[1] = N24 & calc_status_i[86];
  assign N24 = calc_status_i[229] & rs2_match_vector[1];
  assign frs1_data_haz_v[1] = N25 & N26;
  assign N25 = calc_status_i[235] & rs1_match_vector[1];
  assign N26 = calc_status_i[85] | calc_status_i[84];
  assign frs2_data_haz_v[1] = N27 & N28;
  assign N27 = calc_status_i[228] & rs2_match_vector[1];
  assign N28 = calc_status_i[85] | calc_status_i[84];
  assign frs1_data_haz_v[2] = N29 & calc_status_i[94];
  assign N29 = calc_status_i[235] & rs1_match_vector[2];
  assign frs2_data_haz_v[2] = N30 & calc_status_i[94];
  assign N30 = calc_status_i[228] & rs2_match_vector[2];
  assign data_haz_v = N36 | N38;
  assign N36 = N33 | N35;
  assign N33 = N31 | N32;
  assign N31 = irs1_data_haz_v[1] | irs1_data_haz_v[0];
  assign N32 = irs2_data_haz_v[1] | irs2_data_haz_v[0];
  assign N35 = N34 | frs1_data_haz_v[0];
  assign N34 = frs1_data_haz_v[2] | frs1_data_haz_v[1];
  assign N38 = N37 | frs2_data_haz_v[0];
  assign N37 = frs2_data_haz_v[2] | frs2_data_haz_v[1];
  assign struct_haz_v = ~mmu_cmd_ready_i;
  assign mispredict_v = calc_status_i[301] & N6;
  assign chk_dispatch_v_o = ~N39;
  assign N39 = data_haz_v | struct_haz_v;
  assign chk_poison_isd_o = N42 | calc_status_i[1];
  assign N42 = N41 | calc_status_i[2];
  assign N41 = N40 | calc_status_i[3];
  assign N40 = reset_i | mispredict_v;
  assign chk_poison_ex_o = N44 | calc_status_i[1];
  assign N44 = N43 | calc_status_i[2];
  assign N43 = reset_i | calc_status_i[3];

endmodule



module bsg_dff_reset_en_width_p8
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;
  reg [7:0] data_o;
  assign N3 = (N0)? 1'b1 : 
              (N13)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = reset_i;
  assign { N11, N10, N9, N8, N7, N6, N5, N4 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                (N13)? data_i : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N12 = ~reset_i;
  assign N13 = en_i & N12;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[7:0] } <= { N11, N10, N9, N8, N7, N6, N5, N4 };
    end 
  end


endmodule



module bp_be_scheduler_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
(
  clk_i,
  reset_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_o,
  issue_pkt_o,
  issue_pkt_v_o,
  issue_pkt_ready_i
);

  input [133:0] fe_queue_i;
  output [220:0] issue_pkt_o;
  input clk_i;
  input reset_i;
  input fe_queue_v_i;
  input issue_pkt_ready_i;
  output fe_queue_ready_o;
  output issue_pkt_v_o;
  wire [220:0] issue_pkt_o;
  wire fe_queue_ready_o,issue_pkt_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  n_0_net_,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,
  N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298;
  wire [7:0] itag_r,itag_n;
  assign issue_pkt_o[74] = 1'b0;
  assign issue_pkt_o[75] = 1'b0;
  assign issue_pkt_o[212] = fe_queue_i[132];
  assign issue_pkt_o[109] = fe_queue_i[68];
  assign issue_pkt_o[108] = fe_queue_i[67];
  assign issue_pkt_o[107] = fe_queue_i[66];
  assign issue_pkt_o[106] = fe_queue_i[65];
  assign issue_pkt_o[105] = fe_queue_i[64];
  assign issue_pkt_o[104] = fe_queue_i[63];
  assign issue_pkt_o[103] = fe_queue_i[62];
  assign issue_pkt_o[102] = fe_queue_i[61];
  assign issue_pkt_o[101] = fe_queue_i[60];
  assign issue_pkt_o[100] = fe_queue_i[59];
  assign issue_pkt_o[99] = fe_queue_i[58];
  assign issue_pkt_o[98] = fe_queue_i[57];
  assign issue_pkt_o[97] = fe_queue_i[56];
  assign issue_pkt_o[96] = fe_queue_i[55];
  assign issue_pkt_o[95] = fe_queue_i[54];
  assign issue_pkt_o[94] = fe_queue_i[53];
  assign issue_pkt_o[93] = fe_queue_i[52];
  assign issue_pkt_o[92] = fe_queue_i[51];
  assign issue_pkt_o[91] = fe_queue_i[50];
  assign issue_pkt_o[90] = fe_queue_i[49];
  assign issue_pkt_o[89] = fe_queue_i[48];
  assign issue_pkt_o[88] = fe_queue_i[47];
  assign issue_pkt_o[87] = fe_queue_i[46];
  assign issue_pkt_o[86] = fe_queue_i[45];
  assign issue_pkt_o[85] = fe_queue_i[44];
  assign issue_pkt_o[84] = fe_queue_i[43];
  assign issue_pkt_o[83] = fe_queue_i[42];
  assign issue_pkt_o[82] = fe_queue_i[41];
  assign issue_pkt_o[81] = fe_queue_i[40];
  assign issue_pkt_o[80] = fe_queue_i[39];
  assign issue_pkt_o[79] = fe_queue_i[38];
  assign issue_pkt_o[78] = fe_queue_i[37];

  bsg_dff_reset_en_width_p8
  itag_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(n_0_net_),
    .data_i(itag_n),
    .data_o(itag_r)
  );

  assign N15 = fe_queue_i[38] & fe_queue_i[37];
  assign N20 = fe_queue_i[43] | N17;
  assign N21 = N18 | fe_queue_i[40];
  assign N22 = N20 | N21;
  assign N23 = N22 | N19;
  assign N24 = fe_queue_i[43] | fe_queue_i[42];
  assign N25 = N18 | fe_queue_i[40];
  assign N26 = N24 | N25;
  assign N27 = N26 | N19;
  assign N30 = N28 | N17;
  assign N31 = fe_queue_i[41] | N29;
  assign N32 = N30 | N31;
  assign N33 = N32 | N19;
  assign N35 = N28 | N17;
  assign N36 = fe_queue_i[41] | fe_queue_i[40];
  assign N37 = N35 | N36;
  assign N38 = N37 | N19;
  assign N39 = N28 & N17;
  assign N40 = N18 & N29;
  assign N41 = N39 & N40;
  assign N42 = N41 & N19;
  assign N43 = fe_queue_i[43] | fe_queue_i[42];
  assign N44 = N18 | fe_queue_i[40];
  assign N45 = N43 | N44;
  assign N46 = N45 | fe_queue_i[39];
  assign N47 = fe_queue_i[43] | fe_queue_i[42];
  assign N48 = N18 | N29;
  assign N49 = N47 | N48;
  assign N50 = N49 | fe_queue_i[39];
  assign N52 = N28 | N17;
  assign N53 = fe_queue_i[41] | fe_queue_i[40];
  assign N54 = N52 | N53;
  assign N55 = N54 | fe_queue_i[39];
  assign N56 = fe_queue_i[43] | N17;
  assign N57 = fe_queue_i[41] | fe_queue_i[40];
  assign N58 = N56 | N57;
  assign N59 = N58 | fe_queue_i[39];
  assign N60 = fe_queue_i[43] | N17;
  assign N61 = N18 | fe_queue_i[40];
  assign N62 = N60 | N61;
  assign N63 = N62 | fe_queue_i[39];
  assign N64 = fe_queue_i[43] | N17;
  assign N65 = N18 | N29;
  assign N66 = N64 | N65;
  assign N67 = N66 | fe_queue_i[39];
  assign N69 = fe_queue_i[43] & fe_queue_i[41];
  assign N70 = fe_queue_i[41] & fe_queue_i[40];
  assign N71 = N70 & fe_queue_i[39];
  assign N72 = N28 & N18;
  assign N73 = N72 & fe_queue_i[39];
  assign N74 = N17 & N18;
  assign N75 = N74 & fe_queue_i[39];
  assign N76 = N18 & fe_queue_i[40];
  assign N77 = N76 & N19;
  assign N78 = fe_queue_i[43] & N17;
  assign N83 = fe_queue_i[38] & fe_queue_i[37];
  assign N85 = fe_queue_i[43] | N17;
  assign N86 = N18 | fe_queue_i[40];
  assign N87 = N85 | N86;
  assign N88 = N87 | N19;
  assign N89 = fe_queue_i[43] | fe_queue_i[42];
  assign N90 = N18 | fe_queue_i[40];
  assign N91 = N89 | N90;
  assign N92 = N91 | N19;
  assign N94 = N28 | N17;
  assign N95 = fe_queue_i[41] | N29;
  assign N96 = N94 | N95;
  assign N97 = N96 | N19;
  assign N99 = N28 | N17;
  assign N100 = fe_queue_i[41] | fe_queue_i[40];
  assign N101 = N99 | N100;
  assign N102 = N101 | fe_queue_i[39];
  assign N104 = fe_queue_i[43] | N17;
  assign N105 = fe_queue_i[41] | fe_queue_i[40];
  assign N106 = N104 | N105;
  assign N107 = N106 | fe_queue_i[39];
  assign N109 = N28 | N17;
  assign N110 = fe_queue_i[41] | fe_queue_i[40];
  assign N111 = N109 | N110;
  assign N112 = N111 | N19;
  assign N113 = N28 & N17;
  assign N114 = N18 & N29;
  assign N115 = N113 & N114;
  assign N116 = N115 & N19;
  assign N117 = fe_queue_i[43] | fe_queue_i[42];
  assign N118 = N18 | fe_queue_i[40];
  assign N119 = N117 | N118;
  assign N120 = N119 | fe_queue_i[39];
  assign N121 = fe_queue_i[43] | fe_queue_i[42];
  assign N122 = N18 | N29;
  assign N123 = N121 | N122;
  assign N124 = N123 | fe_queue_i[39];
  assign N126 = fe_queue_i[41] & fe_queue_i[40];
  assign N127 = N126 & fe_queue_i[39];
  assign N128 = N28 & N18;
  assign N129 = N128 & fe_queue_i[39];
  assign N130 = N17 & N18;
  assign N131 = N130 & fe_queue_i[39];
  assign N132 = fe_queue_i[43] & fe_queue_i[41];
  assign N133 = fe_queue_i[42] & fe_queue_i[41];
  assign N134 = N133 & N19;
  assign N135 = N18 & fe_queue_i[40];
  assign N136 = N135 & N19;
  assign N137 = fe_queue_i[43] & N17;
  assign N138 = N137 & N19;
  assign itag_n = itag_r + 1'b1;
  assign N80 = (N0)? 1'b0 : 
               (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N34;
  assign N1 = N51;
  assign N2 = N68;
  assign N3 = N79;
  assign { N82, N81 } = (N4)? { N80, N68 } : 
                        (N16)? { 1'b0, 1'b0 } : 1'b0;
  assign N4 = N15;
  assign { N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140 } = (N5)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:49], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N6)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[56:49], fe_queue_i[57:57], fe_queue_i[67:58], 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N7)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[44:44], fe_queue_i[67:62], fe_queue_i[48:45], 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N8)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:62], fe_queue_i[48:44] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:57] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N93;
  assign N6 = N98;
  assign N7 = N103;
  assign N8 = N108;
  assign N9 = N125;
  assign N10 = N139;
  assign { N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204 } = (N11)? { N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = N83;
  assign { issue_pkt_o[220:213], issue_pkt_o[211:149], issue_pkt_o[147:110] } = (N12)? { itag_r, fe_queue_i[131:69], 1'b0, 1'b0, fe_queue_i[36:1] } : 
                                                                                (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:75], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = N14;
  assign N13 = issue_pkt_o[148];
  assign { issue_pkt_o[77:76], issue_pkt_o[73:0] } = (N12)? { N82, N81, fe_queue_i[56:52], fe_queue_i[61:57], N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204 } : 
                                                     (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign fe_queue_ready_o = fe_queue_v_i & issue_pkt_ready_i;
  assign issue_pkt_v_o = fe_queue_v_i & issue_pkt_ready_i;
  assign n_0_net_ = issue_pkt_ready_i & issue_pkt_v_o;
  assign N14 = ~fe_queue_i[133];
  assign issue_pkt_o[148] = fe_queue_i[133];
  assign N16 = ~N15;
  assign N17 = ~fe_queue_i[42];
  assign N18 = ~fe_queue_i[41];
  assign N19 = ~fe_queue_i[39];
  assign N28 = ~fe_queue_i[43];
  assign N29 = ~fe_queue_i[40];
  assign N34 = N270 | N271;
  assign N270 = N268 | N269;
  assign N268 = ~N23;
  assign N269 = ~N27;
  assign N271 = ~N33;
  assign N51 = N275 | N276;
  assign N275 = N273 | N274;
  assign N273 = N272 | N42;
  assign N272 = ~N38;
  assign N274 = ~N46;
  assign N276 = ~N50;
  assign N68 = N281 | N282;
  assign N281 = N279 | N280;
  assign N279 = N277 | N278;
  assign N277 = ~N55;
  assign N278 = ~N59;
  assign N280 = ~N63;
  assign N282 = ~N67;
  assign N79 = N69 | N286;
  assign N286 = N71 | N285;
  assign N285 = N73 | N284;
  assign N284 = N75 | N283;
  assign N283 = N77 | N78;
  assign N84 = ~N83;
  assign N93 = N287 | N288;
  assign N287 = ~N88;
  assign N288 = ~N92;
  assign N98 = ~N97;
  assign N103 = ~N102;
  assign N108 = ~N107;
  assign N125 = N292 | N293;
  assign N292 = N290 | N291;
  assign N290 = N289 | N116;
  assign N289 = ~N112;
  assign N291 = ~N120;
  assign N293 = ~N124;
  assign N139 = N127 | N298;
  assign N298 = N129 | N297;
  assign N297 = N131 | N296;
  assign N296 = N132 | N295;
  assign N295 = N134 | N294;
  assign N294 = N136 | N138;

endmodule



module bp_be_checker_top_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
(
  clk_i,
  reset_i,
  fe_cmd_o,
  fe_cmd_v_o,
  fe_cmd_ready_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_o,
  chk_roll_fe_o,
  chk_flush_fe_o,
  chk_dequeue_fe_o,
  issue_pkt_o,
  issue_pkt_v_o,
  issue_pkt_ready_i,
  calc_status_i,
  mmu_cmd_ready_i,
  chk_dispatch_v_o,
  chk_roll_o,
  chk_poison_isd_o,
  chk_poison_ex_o
);

  output [108:0] fe_cmd_o;
  input [133:0] fe_queue_i;
  output [220:0] issue_pkt_o;
  input [301:0] calc_status_i;
  input clk_i;
  input reset_i;
  input fe_cmd_ready_i;
  input fe_queue_v_i;
  input issue_pkt_ready_i;
  input mmu_cmd_ready_i;
  output fe_cmd_v_o;
  output fe_queue_ready_o;
  output chk_roll_fe_o;
  output chk_flush_fe_o;
  output chk_dequeue_fe_o;
  output issue_pkt_v_o;
  output chk_dispatch_v_o;
  output chk_roll_o;
  output chk_poison_isd_o;
  output chk_poison_ex_o;
  wire [108:0] fe_cmd_o;
  wire [220:0] issue_pkt_o;
  wire fe_cmd_v_o,fe_queue_ready_o,chk_roll_fe_o,chk_flush_fe_o,chk_dequeue_fe_o,
  issue_pkt_v_o,chk_dispatch_v_o,chk_roll_o,chk_poison_isd_o,chk_poison_ex_o;
  wire [63:0] expected_npc;

  bp_be_director_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
  director
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .calc_status_i(calc_status_i),
    .expected_npc_o(expected_npc),
    .fe_cmd_o(fe_cmd_o),
    .fe_cmd_v_o(fe_cmd_v_o),
    .fe_cmd_ready_i(fe_cmd_ready_i),
    .chk_flush_fe_o(chk_flush_fe_o),
    .chk_dequeue_fe_o(chk_dequeue_fe_o),
    .chk_roll_fe_o(chk_roll_fe_o)
  );


  bp_be_detector_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
  detector
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .calc_status_i(calc_status_i),
    .expected_npc_i(expected_npc),
    .mmu_cmd_ready_i(mmu_cmd_ready_i),
    .chk_dispatch_v_o(chk_dispatch_v_o),
    .chk_roll_o(chk_roll_o),
    .chk_poison_isd_o(chk_poison_isd_o),
    .chk_poison_ex_o(chk_poison_ex_o)
  );


  bp_be_scheduler_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
  scheduler
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fe_queue_i(fe_queue_i),
    .fe_queue_v_i(fe_queue_v_i),
    .fe_queue_ready_o(fe_queue_ready_o),
    .issue_pkt_o(issue_pkt_o),
    .issue_pkt_v_o(issue_pkt_v_o),
    .issue_pkt_ready_i(issue_pkt_ready_i)
  );


endmodule



module bsg_mem_2r1w_sync_synth_width_p64_els_p32_read_write_same_addr_p1_harden_p0
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r0_v_i,
  r0_addr_i,
  r0_data_o,
  r1_v_i,
  r1_addr_i,
  r1_data_o
);

  input [4:0] w_addr_i;
  input [63:0] w_data_i;
  input [4:0] r0_addr_i;
  output [63:0] r0_data_o;
  input [4:0] r1_addr_i;
  output [63:0] r1_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r0_v_i;
  input r1_v_i;
  wire [63:0] r0_data_o,r1_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221;
  reg [4:0] r0_addr_r,r1_addr_r;
  reg [2047:0] mem;
  assign r0_data_o[63] = (N43)? mem[63] : 
                         (N45)? mem[127] : 
                         (N47)? mem[191] : 
                         (N49)? mem[255] : 
                         (N51)? mem[319] : 
                         (N53)? mem[383] : 
                         (N55)? mem[447] : 
                         (N57)? mem[511] : 
                         (N59)? mem[575] : 
                         (N61)? mem[639] : 
                         (N63)? mem[703] : 
                         (N65)? mem[767] : 
                         (N67)? mem[831] : 
                         (N69)? mem[895] : 
                         (N71)? mem[959] : 
                         (N73)? mem[1023] : 
                         (N44)? mem[1087] : 
                         (N46)? mem[1151] : 
                         (N48)? mem[1215] : 
                         (N50)? mem[1279] : 
                         (N52)? mem[1343] : 
                         (N54)? mem[1407] : 
                         (N56)? mem[1471] : 
                         (N58)? mem[1535] : 
                         (N60)? mem[1599] : 
                         (N62)? mem[1663] : 
                         (N64)? mem[1727] : 
                         (N66)? mem[1791] : 
                         (N68)? mem[1855] : 
                         (N70)? mem[1919] : 
                         (N72)? mem[1983] : 
                         (N74)? mem[2047] : 1'b0;
  assign r0_data_o[62] = (N43)? mem[62] : 
                         (N45)? mem[126] : 
                         (N47)? mem[190] : 
                         (N49)? mem[254] : 
                         (N51)? mem[318] : 
                         (N53)? mem[382] : 
                         (N55)? mem[446] : 
                         (N57)? mem[510] : 
                         (N59)? mem[574] : 
                         (N61)? mem[638] : 
                         (N63)? mem[702] : 
                         (N65)? mem[766] : 
                         (N67)? mem[830] : 
                         (N69)? mem[894] : 
                         (N71)? mem[958] : 
                         (N73)? mem[1022] : 
                         (N44)? mem[1086] : 
                         (N46)? mem[1150] : 
                         (N48)? mem[1214] : 
                         (N50)? mem[1278] : 
                         (N52)? mem[1342] : 
                         (N54)? mem[1406] : 
                         (N56)? mem[1470] : 
                         (N58)? mem[1534] : 
                         (N60)? mem[1598] : 
                         (N62)? mem[1662] : 
                         (N64)? mem[1726] : 
                         (N66)? mem[1790] : 
                         (N68)? mem[1854] : 
                         (N70)? mem[1918] : 
                         (N72)? mem[1982] : 
                         (N74)? mem[2046] : 1'b0;
  assign r0_data_o[61] = (N43)? mem[61] : 
                         (N45)? mem[125] : 
                         (N47)? mem[189] : 
                         (N49)? mem[253] : 
                         (N51)? mem[317] : 
                         (N53)? mem[381] : 
                         (N55)? mem[445] : 
                         (N57)? mem[509] : 
                         (N59)? mem[573] : 
                         (N61)? mem[637] : 
                         (N63)? mem[701] : 
                         (N65)? mem[765] : 
                         (N67)? mem[829] : 
                         (N69)? mem[893] : 
                         (N71)? mem[957] : 
                         (N73)? mem[1021] : 
                         (N44)? mem[1085] : 
                         (N46)? mem[1149] : 
                         (N48)? mem[1213] : 
                         (N50)? mem[1277] : 
                         (N52)? mem[1341] : 
                         (N54)? mem[1405] : 
                         (N56)? mem[1469] : 
                         (N58)? mem[1533] : 
                         (N60)? mem[1597] : 
                         (N62)? mem[1661] : 
                         (N64)? mem[1725] : 
                         (N66)? mem[1789] : 
                         (N68)? mem[1853] : 
                         (N70)? mem[1917] : 
                         (N72)? mem[1981] : 
                         (N74)? mem[2045] : 1'b0;
  assign r0_data_o[60] = (N43)? mem[60] : 
                         (N45)? mem[124] : 
                         (N47)? mem[188] : 
                         (N49)? mem[252] : 
                         (N51)? mem[316] : 
                         (N53)? mem[380] : 
                         (N55)? mem[444] : 
                         (N57)? mem[508] : 
                         (N59)? mem[572] : 
                         (N61)? mem[636] : 
                         (N63)? mem[700] : 
                         (N65)? mem[764] : 
                         (N67)? mem[828] : 
                         (N69)? mem[892] : 
                         (N71)? mem[956] : 
                         (N73)? mem[1020] : 
                         (N44)? mem[1084] : 
                         (N46)? mem[1148] : 
                         (N48)? mem[1212] : 
                         (N50)? mem[1276] : 
                         (N52)? mem[1340] : 
                         (N54)? mem[1404] : 
                         (N56)? mem[1468] : 
                         (N58)? mem[1532] : 
                         (N60)? mem[1596] : 
                         (N62)? mem[1660] : 
                         (N64)? mem[1724] : 
                         (N66)? mem[1788] : 
                         (N68)? mem[1852] : 
                         (N70)? mem[1916] : 
                         (N72)? mem[1980] : 
                         (N74)? mem[2044] : 1'b0;
  assign r0_data_o[59] = (N43)? mem[59] : 
                         (N45)? mem[123] : 
                         (N47)? mem[187] : 
                         (N49)? mem[251] : 
                         (N51)? mem[315] : 
                         (N53)? mem[379] : 
                         (N55)? mem[443] : 
                         (N57)? mem[507] : 
                         (N59)? mem[571] : 
                         (N61)? mem[635] : 
                         (N63)? mem[699] : 
                         (N65)? mem[763] : 
                         (N67)? mem[827] : 
                         (N69)? mem[891] : 
                         (N71)? mem[955] : 
                         (N73)? mem[1019] : 
                         (N44)? mem[1083] : 
                         (N46)? mem[1147] : 
                         (N48)? mem[1211] : 
                         (N50)? mem[1275] : 
                         (N52)? mem[1339] : 
                         (N54)? mem[1403] : 
                         (N56)? mem[1467] : 
                         (N58)? mem[1531] : 
                         (N60)? mem[1595] : 
                         (N62)? mem[1659] : 
                         (N64)? mem[1723] : 
                         (N66)? mem[1787] : 
                         (N68)? mem[1851] : 
                         (N70)? mem[1915] : 
                         (N72)? mem[1979] : 
                         (N74)? mem[2043] : 1'b0;
  assign r0_data_o[58] = (N43)? mem[58] : 
                         (N45)? mem[122] : 
                         (N47)? mem[186] : 
                         (N49)? mem[250] : 
                         (N51)? mem[314] : 
                         (N53)? mem[378] : 
                         (N55)? mem[442] : 
                         (N57)? mem[506] : 
                         (N59)? mem[570] : 
                         (N61)? mem[634] : 
                         (N63)? mem[698] : 
                         (N65)? mem[762] : 
                         (N67)? mem[826] : 
                         (N69)? mem[890] : 
                         (N71)? mem[954] : 
                         (N73)? mem[1018] : 
                         (N44)? mem[1082] : 
                         (N46)? mem[1146] : 
                         (N48)? mem[1210] : 
                         (N50)? mem[1274] : 
                         (N52)? mem[1338] : 
                         (N54)? mem[1402] : 
                         (N56)? mem[1466] : 
                         (N58)? mem[1530] : 
                         (N60)? mem[1594] : 
                         (N62)? mem[1658] : 
                         (N64)? mem[1722] : 
                         (N66)? mem[1786] : 
                         (N68)? mem[1850] : 
                         (N70)? mem[1914] : 
                         (N72)? mem[1978] : 
                         (N74)? mem[2042] : 1'b0;
  assign r0_data_o[57] = (N43)? mem[57] : 
                         (N45)? mem[121] : 
                         (N47)? mem[185] : 
                         (N49)? mem[249] : 
                         (N51)? mem[313] : 
                         (N53)? mem[377] : 
                         (N55)? mem[441] : 
                         (N57)? mem[505] : 
                         (N59)? mem[569] : 
                         (N61)? mem[633] : 
                         (N63)? mem[697] : 
                         (N65)? mem[761] : 
                         (N67)? mem[825] : 
                         (N69)? mem[889] : 
                         (N71)? mem[953] : 
                         (N73)? mem[1017] : 
                         (N44)? mem[1081] : 
                         (N46)? mem[1145] : 
                         (N48)? mem[1209] : 
                         (N50)? mem[1273] : 
                         (N52)? mem[1337] : 
                         (N54)? mem[1401] : 
                         (N56)? mem[1465] : 
                         (N58)? mem[1529] : 
                         (N60)? mem[1593] : 
                         (N62)? mem[1657] : 
                         (N64)? mem[1721] : 
                         (N66)? mem[1785] : 
                         (N68)? mem[1849] : 
                         (N70)? mem[1913] : 
                         (N72)? mem[1977] : 
                         (N74)? mem[2041] : 1'b0;
  assign r0_data_o[56] = (N43)? mem[56] : 
                         (N45)? mem[120] : 
                         (N47)? mem[184] : 
                         (N49)? mem[248] : 
                         (N51)? mem[312] : 
                         (N53)? mem[376] : 
                         (N55)? mem[440] : 
                         (N57)? mem[504] : 
                         (N59)? mem[568] : 
                         (N61)? mem[632] : 
                         (N63)? mem[696] : 
                         (N65)? mem[760] : 
                         (N67)? mem[824] : 
                         (N69)? mem[888] : 
                         (N71)? mem[952] : 
                         (N73)? mem[1016] : 
                         (N44)? mem[1080] : 
                         (N46)? mem[1144] : 
                         (N48)? mem[1208] : 
                         (N50)? mem[1272] : 
                         (N52)? mem[1336] : 
                         (N54)? mem[1400] : 
                         (N56)? mem[1464] : 
                         (N58)? mem[1528] : 
                         (N60)? mem[1592] : 
                         (N62)? mem[1656] : 
                         (N64)? mem[1720] : 
                         (N66)? mem[1784] : 
                         (N68)? mem[1848] : 
                         (N70)? mem[1912] : 
                         (N72)? mem[1976] : 
                         (N74)? mem[2040] : 1'b0;
  assign r0_data_o[55] = (N43)? mem[55] : 
                         (N45)? mem[119] : 
                         (N47)? mem[183] : 
                         (N49)? mem[247] : 
                         (N51)? mem[311] : 
                         (N53)? mem[375] : 
                         (N55)? mem[439] : 
                         (N57)? mem[503] : 
                         (N59)? mem[567] : 
                         (N61)? mem[631] : 
                         (N63)? mem[695] : 
                         (N65)? mem[759] : 
                         (N67)? mem[823] : 
                         (N69)? mem[887] : 
                         (N71)? mem[951] : 
                         (N73)? mem[1015] : 
                         (N44)? mem[1079] : 
                         (N46)? mem[1143] : 
                         (N48)? mem[1207] : 
                         (N50)? mem[1271] : 
                         (N52)? mem[1335] : 
                         (N54)? mem[1399] : 
                         (N56)? mem[1463] : 
                         (N58)? mem[1527] : 
                         (N60)? mem[1591] : 
                         (N62)? mem[1655] : 
                         (N64)? mem[1719] : 
                         (N66)? mem[1783] : 
                         (N68)? mem[1847] : 
                         (N70)? mem[1911] : 
                         (N72)? mem[1975] : 
                         (N74)? mem[2039] : 1'b0;
  assign r0_data_o[54] = (N43)? mem[54] : 
                         (N45)? mem[118] : 
                         (N47)? mem[182] : 
                         (N49)? mem[246] : 
                         (N51)? mem[310] : 
                         (N53)? mem[374] : 
                         (N55)? mem[438] : 
                         (N57)? mem[502] : 
                         (N59)? mem[566] : 
                         (N61)? mem[630] : 
                         (N63)? mem[694] : 
                         (N65)? mem[758] : 
                         (N67)? mem[822] : 
                         (N69)? mem[886] : 
                         (N71)? mem[950] : 
                         (N73)? mem[1014] : 
                         (N44)? mem[1078] : 
                         (N46)? mem[1142] : 
                         (N48)? mem[1206] : 
                         (N50)? mem[1270] : 
                         (N52)? mem[1334] : 
                         (N54)? mem[1398] : 
                         (N56)? mem[1462] : 
                         (N58)? mem[1526] : 
                         (N60)? mem[1590] : 
                         (N62)? mem[1654] : 
                         (N64)? mem[1718] : 
                         (N66)? mem[1782] : 
                         (N68)? mem[1846] : 
                         (N70)? mem[1910] : 
                         (N72)? mem[1974] : 
                         (N74)? mem[2038] : 1'b0;
  assign r0_data_o[53] = (N43)? mem[53] : 
                         (N45)? mem[117] : 
                         (N47)? mem[181] : 
                         (N49)? mem[245] : 
                         (N51)? mem[309] : 
                         (N53)? mem[373] : 
                         (N55)? mem[437] : 
                         (N57)? mem[501] : 
                         (N59)? mem[565] : 
                         (N61)? mem[629] : 
                         (N63)? mem[693] : 
                         (N65)? mem[757] : 
                         (N67)? mem[821] : 
                         (N69)? mem[885] : 
                         (N71)? mem[949] : 
                         (N73)? mem[1013] : 
                         (N44)? mem[1077] : 
                         (N46)? mem[1141] : 
                         (N48)? mem[1205] : 
                         (N50)? mem[1269] : 
                         (N52)? mem[1333] : 
                         (N54)? mem[1397] : 
                         (N56)? mem[1461] : 
                         (N58)? mem[1525] : 
                         (N60)? mem[1589] : 
                         (N62)? mem[1653] : 
                         (N64)? mem[1717] : 
                         (N66)? mem[1781] : 
                         (N68)? mem[1845] : 
                         (N70)? mem[1909] : 
                         (N72)? mem[1973] : 
                         (N74)? mem[2037] : 1'b0;
  assign r0_data_o[52] = (N43)? mem[52] : 
                         (N45)? mem[116] : 
                         (N47)? mem[180] : 
                         (N49)? mem[244] : 
                         (N51)? mem[308] : 
                         (N53)? mem[372] : 
                         (N55)? mem[436] : 
                         (N57)? mem[500] : 
                         (N59)? mem[564] : 
                         (N61)? mem[628] : 
                         (N63)? mem[692] : 
                         (N65)? mem[756] : 
                         (N67)? mem[820] : 
                         (N69)? mem[884] : 
                         (N71)? mem[948] : 
                         (N73)? mem[1012] : 
                         (N44)? mem[1076] : 
                         (N46)? mem[1140] : 
                         (N48)? mem[1204] : 
                         (N50)? mem[1268] : 
                         (N52)? mem[1332] : 
                         (N54)? mem[1396] : 
                         (N56)? mem[1460] : 
                         (N58)? mem[1524] : 
                         (N60)? mem[1588] : 
                         (N62)? mem[1652] : 
                         (N64)? mem[1716] : 
                         (N66)? mem[1780] : 
                         (N68)? mem[1844] : 
                         (N70)? mem[1908] : 
                         (N72)? mem[1972] : 
                         (N74)? mem[2036] : 1'b0;
  assign r0_data_o[51] = (N43)? mem[51] : 
                         (N45)? mem[115] : 
                         (N47)? mem[179] : 
                         (N49)? mem[243] : 
                         (N51)? mem[307] : 
                         (N53)? mem[371] : 
                         (N55)? mem[435] : 
                         (N57)? mem[499] : 
                         (N59)? mem[563] : 
                         (N61)? mem[627] : 
                         (N63)? mem[691] : 
                         (N65)? mem[755] : 
                         (N67)? mem[819] : 
                         (N69)? mem[883] : 
                         (N71)? mem[947] : 
                         (N73)? mem[1011] : 
                         (N44)? mem[1075] : 
                         (N46)? mem[1139] : 
                         (N48)? mem[1203] : 
                         (N50)? mem[1267] : 
                         (N52)? mem[1331] : 
                         (N54)? mem[1395] : 
                         (N56)? mem[1459] : 
                         (N58)? mem[1523] : 
                         (N60)? mem[1587] : 
                         (N62)? mem[1651] : 
                         (N64)? mem[1715] : 
                         (N66)? mem[1779] : 
                         (N68)? mem[1843] : 
                         (N70)? mem[1907] : 
                         (N72)? mem[1971] : 
                         (N74)? mem[2035] : 1'b0;
  assign r0_data_o[50] = (N43)? mem[50] : 
                         (N45)? mem[114] : 
                         (N47)? mem[178] : 
                         (N49)? mem[242] : 
                         (N51)? mem[306] : 
                         (N53)? mem[370] : 
                         (N55)? mem[434] : 
                         (N57)? mem[498] : 
                         (N59)? mem[562] : 
                         (N61)? mem[626] : 
                         (N63)? mem[690] : 
                         (N65)? mem[754] : 
                         (N67)? mem[818] : 
                         (N69)? mem[882] : 
                         (N71)? mem[946] : 
                         (N73)? mem[1010] : 
                         (N44)? mem[1074] : 
                         (N46)? mem[1138] : 
                         (N48)? mem[1202] : 
                         (N50)? mem[1266] : 
                         (N52)? mem[1330] : 
                         (N54)? mem[1394] : 
                         (N56)? mem[1458] : 
                         (N58)? mem[1522] : 
                         (N60)? mem[1586] : 
                         (N62)? mem[1650] : 
                         (N64)? mem[1714] : 
                         (N66)? mem[1778] : 
                         (N68)? mem[1842] : 
                         (N70)? mem[1906] : 
                         (N72)? mem[1970] : 
                         (N74)? mem[2034] : 1'b0;
  assign r0_data_o[49] = (N43)? mem[49] : 
                         (N45)? mem[113] : 
                         (N47)? mem[177] : 
                         (N49)? mem[241] : 
                         (N51)? mem[305] : 
                         (N53)? mem[369] : 
                         (N55)? mem[433] : 
                         (N57)? mem[497] : 
                         (N59)? mem[561] : 
                         (N61)? mem[625] : 
                         (N63)? mem[689] : 
                         (N65)? mem[753] : 
                         (N67)? mem[817] : 
                         (N69)? mem[881] : 
                         (N71)? mem[945] : 
                         (N73)? mem[1009] : 
                         (N44)? mem[1073] : 
                         (N46)? mem[1137] : 
                         (N48)? mem[1201] : 
                         (N50)? mem[1265] : 
                         (N52)? mem[1329] : 
                         (N54)? mem[1393] : 
                         (N56)? mem[1457] : 
                         (N58)? mem[1521] : 
                         (N60)? mem[1585] : 
                         (N62)? mem[1649] : 
                         (N64)? mem[1713] : 
                         (N66)? mem[1777] : 
                         (N68)? mem[1841] : 
                         (N70)? mem[1905] : 
                         (N72)? mem[1969] : 
                         (N74)? mem[2033] : 1'b0;
  assign r0_data_o[48] = (N43)? mem[48] : 
                         (N45)? mem[112] : 
                         (N47)? mem[176] : 
                         (N49)? mem[240] : 
                         (N51)? mem[304] : 
                         (N53)? mem[368] : 
                         (N55)? mem[432] : 
                         (N57)? mem[496] : 
                         (N59)? mem[560] : 
                         (N61)? mem[624] : 
                         (N63)? mem[688] : 
                         (N65)? mem[752] : 
                         (N67)? mem[816] : 
                         (N69)? mem[880] : 
                         (N71)? mem[944] : 
                         (N73)? mem[1008] : 
                         (N44)? mem[1072] : 
                         (N46)? mem[1136] : 
                         (N48)? mem[1200] : 
                         (N50)? mem[1264] : 
                         (N52)? mem[1328] : 
                         (N54)? mem[1392] : 
                         (N56)? mem[1456] : 
                         (N58)? mem[1520] : 
                         (N60)? mem[1584] : 
                         (N62)? mem[1648] : 
                         (N64)? mem[1712] : 
                         (N66)? mem[1776] : 
                         (N68)? mem[1840] : 
                         (N70)? mem[1904] : 
                         (N72)? mem[1968] : 
                         (N74)? mem[2032] : 1'b0;
  assign r0_data_o[47] = (N43)? mem[47] : 
                         (N45)? mem[111] : 
                         (N47)? mem[175] : 
                         (N49)? mem[239] : 
                         (N51)? mem[303] : 
                         (N53)? mem[367] : 
                         (N55)? mem[431] : 
                         (N57)? mem[495] : 
                         (N59)? mem[559] : 
                         (N61)? mem[623] : 
                         (N63)? mem[687] : 
                         (N65)? mem[751] : 
                         (N67)? mem[815] : 
                         (N69)? mem[879] : 
                         (N71)? mem[943] : 
                         (N73)? mem[1007] : 
                         (N44)? mem[1071] : 
                         (N46)? mem[1135] : 
                         (N48)? mem[1199] : 
                         (N50)? mem[1263] : 
                         (N52)? mem[1327] : 
                         (N54)? mem[1391] : 
                         (N56)? mem[1455] : 
                         (N58)? mem[1519] : 
                         (N60)? mem[1583] : 
                         (N62)? mem[1647] : 
                         (N64)? mem[1711] : 
                         (N66)? mem[1775] : 
                         (N68)? mem[1839] : 
                         (N70)? mem[1903] : 
                         (N72)? mem[1967] : 
                         (N74)? mem[2031] : 1'b0;
  assign r0_data_o[46] = (N43)? mem[46] : 
                         (N45)? mem[110] : 
                         (N47)? mem[174] : 
                         (N49)? mem[238] : 
                         (N51)? mem[302] : 
                         (N53)? mem[366] : 
                         (N55)? mem[430] : 
                         (N57)? mem[494] : 
                         (N59)? mem[558] : 
                         (N61)? mem[622] : 
                         (N63)? mem[686] : 
                         (N65)? mem[750] : 
                         (N67)? mem[814] : 
                         (N69)? mem[878] : 
                         (N71)? mem[942] : 
                         (N73)? mem[1006] : 
                         (N44)? mem[1070] : 
                         (N46)? mem[1134] : 
                         (N48)? mem[1198] : 
                         (N50)? mem[1262] : 
                         (N52)? mem[1326] : 
                         (N54)? mem[1390] : 
                         (N56)? mem[1454] : 
                         (N58)? mem[1518] : 
                         (N60)? mem[1582] : 
                         (N62)? mem[1646] : 
                         (N64)? mem[1710] : 
                         (N66)? mem[1774] : 
                         (N68)? mem[1838] : 
                         (N70)? mem[1902] : 
                         (N72)? mem[1966] : 
                         (N74)? mem[2030] : 1'b0;
  assign r0_data_o[45] = (N43)? mem[45] : 
                         (N45)? mem[109] : 
                         (N47)? mem[173] : 
                         (N49)? mem[237] : 
                         (N51)? mem[301] : 
                         (N53)? mem[365] : 
                         (N55)? mem[429] : 
                         (N57)? mem[493] : 
                         (N59)? mem[557] : 
                         (N61)? mem[621] : 
                         (N63)? mem[685] : 
                         (N65)? mem[749] : 
                         (N67)? mem[813] : 
                         (N69)? mem[877] : 
                         (N71)? mem[941] : 
                         (N73)? mem[1005] : 
                         (N44)? mem[1069] : 
                         (N46)? mem[1133] : 
                         (N48)? mem[1197] : 
                         (N50)? mem[1261] : 
                         (N52)? mem[1325] : 
                         (N54)? mem[1389] : 
                         (N56)? mem[1453] : 
                         (N58)? mem[1517] : 
                         (N60)? mem[1581] : 
                         (N62)? mem[1645] : 
                         (N64)? mem[1709] : 
                         (N66)? mem[1773] : 
                         (N68)? mem[1837] : 
                         (N70)? mem[1901] : 
                         (N72)? mem[1965] : 
                         (N74)? mem[2029] : 1'b0;
  assign r0_data_o[44] = (N43)? mem[44] : 
                         (N45)? mem[108] : 
                         (N47)? mem[172] : 
                         (N49)? mem[236] : 
                         (N51)? mem[300] : 
                         (N53)? mem[364] : 
                         (N55)? mem[428] : 
                         (N57)? mem[492] : 
                         (N59)? mem[556] : 
                         (N61)? mem[620] : 
                         (N63)? mem[684] : 
                         (N65)? mem[748] : 
                         (N67)? mem[812] : 
                         (N69)? mem[876] : 
                         (N71)? mem[940] : 
                         (N73)? mem[1004] : 
                         (N44)? mem[1068] : 
                         (N46)? mem[1132] : 
                         (N48)? mem[1196] : 
                         (N50)? mem[1260] : 
                         (N52)? mem[1324] : 
                         (N54)? mem[1388] : 
                         (N56)? mem[1452] : 
                         (N58)? mem[1516] : 
                         (N60)? mem[1580] : 
                         (N62)? mem[1644] : 
                         (N64)? mem[1708] : 
                         (N66)? mem[1772] : 
                         (N68)? mem[1836] : 
                         (N70)? mem[1900] : 
                         (N72)? mem[1964] : 
                         (N74)? mem[2028] : 1'b0;
  assign r0_data_o[43] = (N43)? mem[43] : 
                         (N45)? mem[107] : 
                         (N47)? mem[171] : 
                         (N49)? mem[235] : 
                         (N51)? mem[299] : 
                         (N53)? mem[363] : 
                         (N55)? mem[427] : 
                         (N57)? mem[491] : 
                         (N59)? mem[555] : 
                         (N61)? mem[619] : 
                         (N63)? mem[683] : 
                         (N65)? mem[747] : 
                         (N67)? mem[811] : 
                         (N69)? mem[875] : 
                         (N71)? mem[939] : 
                         (N73)? mem[1003] : 
                         (N44)? mem[1067] : 
                         (N46)? mem[1131] : 
                         (N48)? mem[1195] : 
                         (N50)? mem[1259] : 
                         (N52)? mem[1323] : 
                         (N54)? mem[1387] : 
                         (N56)? mem[1451] : 
                         (N58)? mem[1515] : 
                         (N60)? mem[1579] : 
                         (N62)? mem[1643] : 
                         (N64)? mem[1707] : 
                         (N66)? mem[1771] : 
                         (N68)? mem[1835] : 
                         (N70)? mem[1899] : 
                         (N72)? mem[1963] : 
                         (N74)? mem[2027] : 1'b0;
  assign r0_data_o[42] = (N43)? mem[42] : 
                         (N45)? mem[106] : 
                         (N47)? mem[170] : 
                         (N49)? mem[234] : 
                         (N51)? mem[298] : 
                         (N53)? mem[362] : 
                         (N55)? mem[426] : 
                         (N57)? mem[490] : 
                         (N59)? mem[554] : 
                         (N61)? mem[618] : 
                         (N63)? mem[682] : 
                         (N65)? mem[746] : 
                         (N67)? mem[810] : 
                         (N69)? mem[874] : 
                         (N71)? mem[938] : 
                         (N73)? mem[1002] : 
                         (N44)? mem[1066] : 
                         (N46)? mem[1130] : 
                         (N48)? mem[1194] : 
                         (N50)? mem[1258] : 
                         (N52)? mem[1322] : 
                         (N54)? mem[1386] : 
                         (N56)? mem[1450] : 
                         (N58)? mem[1514] : 
                         (N60)? mem[1578] : 
                         (N62)? mem[1642] : 
                         (N64)? mem[1706] : 
                         (N66)? mem[1770] : 
                         (N68)? mem[1834] : 
                         (N70)? mem[1898] : 
                         (N72)? mem[1962] : 
                         (N74)? mem[2026] : 1'b0;
  assign r0_data_o[41] = (N43)? mem[41] : 
                         (N45)? mem[105] : 
                         (N47)? mem[169] : 
                         (N49)? mem[233] : 
                         (N51)? mem[297] : 
                         (N53)? mem[361] : 
                         (N55)? mem[425] : 
                         (N57)? mem[489] : 
                         (N59)? mem[553] : 
                         (N61)? mem[617] : 
                         (N63)? mem[681] : 
                         (N65)? mem[745] : 
                         (N67)? mem[809] : 
                         (N69)? mem[873] : 
                         (N71)? mem[937] : 
                         (N73)? mem[1001] : 
                         (N44)? mem[1065] : 
                         (N46)? mem[1129] : 
                         (N48)? mem[1193] : 
                         (N50)? mem[1257] : 
                         (N52)? mem[1321] : 
                         (N54)? mem[1385] : 
                         (N56)? mem[1449] : 
                         (N58)? mem[1513] : 
                         (N60)? mem[1577] : 
                         (N62)? mem[1641] : 
                         (N64)? mem[1705] : 
                         (N66)? mem[1769] : 
                         (N68)? mem[1833] : 
                         (N70)? mem[1897] : 
                         (N72)? mem[1961] : 
                         (N74)? mem[2025] : 1'b0;
  assign r0_data_o[40] = (N43)? mem[40] : 
                         (N45)? mem[104] : 
                         (N47)? mem[168] : 
                         (N49)? mem[232] : 
                         (N51)? mem[296] : 
                         (N53)? mem[360] : 
                         (N55)? mem[424] : 
                         (N57)? mem[488] : 
                         (N59)? mem[552] : 
                         (N61)? mem[616] : 
                         (N63)? mem[680] : 
                         (N65)? mem[744] : 
                         (N67)? mem[808] : 
                         (N69)? mem[872] : 
                         (N71)? mem[936] : 
                         (N73)? mem[1000] : 
                         (N44)? mem[1064] : 
                         (N46)? mem[1128] : 
                         (N48)? mem[1192] : 
                         (N50)? mem[1256] : 
                         (N52)? mem[1320] : 
                         (N54)? mem[1384] : 
                         (N56)? mem[1448] : 
                         (N58)? mem[1512] : 
                         (N60)? mem[1576] : 
                         (N62)? mem[1640] : 
                         (N64)? mem[1704] : 
                         (N66)? mem[1768] : 
                         (N68)? mem[1832] : 
                         (N70)? mem[1896] : 
                         (N72)? mem[1960] : 
                         (N74)? mem[2024] : 1'b0;
  assign r0_data_o[39] = (N43)? mem[39] : 
                         (N45)? mem[103] : 
                         (N47)? mem[167] : 
                         (N49)? mem[231] : 
                         (N51)? mem[295] : 
                         (N53)? mem[359] : 
                         (N55)? mem[423] : 
                         (N57)? mem[487] : 
                         (N59)? mem[551] : 
                         (N61)? mem[615] : 
                         (N63)? mem[679] : 
                         (N65)? mem[743] : 
                         (N67)? mem[807] : 
                         (N69)? mem[871] : 
                         (N71)? mem[935] : 
                         (N73)? mem[999] : 
                         (N44)? mem[1063] : 
                         (N46)? mem[1127] : 
                         (N48)? mem[1191] : 
                         (N50)? mem[1255] : 
                         (N52)? mem[1319] : 
                         (N54)? mem[1383] : 
                         (N56)? mem[1447] : 
                         (N58)? mem[1511] : 
                         (N60)? mem[1575] : 
                         (N62)? mem[1639] : 
                         (N64)? mem[1703] : 
                         (N66)? mem[1767] : 
                         (N68)? mem[1831] : 
                         (N70)? mem[1895] : 
                         (N72)? mem[1959] : 
                         (N74)? mem[2023] : 1'b0;
  assign r0_data_o[38] = (N43)? mem[38] : 
                         (N45)? mem[102] : 
                         (N47)? mem[166] : 
                         (N49)? mem[230] : 
                         (N51)? mem[294] : 
                         (N53)? mem[358] : 
                         (N55)? mem[422] : 
                         (N57)? mem[486] : 
                         (N59)? mem[550] : 
                         (N61)? mem[614] : 
                         (N63)? mem[678] : 
                         (N65)? mem[742] : 
                         (N67)? mem[806] : 
                         (N69)? mem[870] : 
                         (N71)? mem[934] : 
                         (N73)? mem[998] : 
                         (N44)? mem[1062] : 
                         (N46)? mem[1126] : 
                         (N48)? mem[1190] : 
                         (N50)? mem[1254] : 
                         (N52)? mem[1318] : 
                         (N54)? mem[1382] : 
                         (N56)? mem[1446] : 
                         (N58)? mem[1510] : 
                         (N60)? mem[1574] : 
                         (N62)? mem[1638] : 
                         (N64)? mem[1702] : 
                         (N66)? mem[1766] : 
                         (N68)? mem[1830] : 
                         (N70)? mem[1894] : 
                         (N72)? mem[1958] : 
                         (N74)? mem[2022] : 1'b0;
  assign r0_data_o[37] = (N43)? mem[37] : 
                         (N45)? mem[101] : 
                         (N47)? mem[165] : 
                         (N49)? mem[229] : 
                         (N51)? mem[293] : 
                         (N53)? mem[357] : 
                         (N55)? mem[421] : 
                         (N57)? mem[485] : 
                         (N59)? mem[549] : 
                         (N61)? mem[613] : 
                         (N63)? mem[677] : 
                         (N65)? mem[741] : 
                         (N67)? mem[805] : 
                         (N69)? mem[869] : 
                         (N71)? mem[933] : 
                         (N73)? mem[997] : 
                         (N44)? mem[1061] : 
                         (N46)? mem[1125] : 
                         (N48)? mem[1189] : 
                         (N50)? mem[1253] : 
                         (N52)? mem[1317] : 
                         (N54)? mem[1381] : 
                         (N56)? mem[1445] : 
                         (N58)? mem[1509] : 
                         (N60)? mem[1573] : 
                         (N62)? mem[1637] : 
                         (N64)? mem[1701] : 
                         (N66)? mem[1765] : 
                         (N68)? mem[1829] : 
                         (N70)? mem[1893] : 
                         (N72)? mem[1957] : 
                         (N74)? mem[2021] : 1'b0;
  assign r0_data_o[36] = (N43)? mem[36] : 
                         (N45)? mem[100] : 
                         (N47)? mem[164] : 
                         (N49)? mem[228] : 
                         (N51)? mem[292] : 
                         (N53)? mem[356] : 
                         (N55)? mem[420] : 
                         (N57)? mem[484] : 
                         (N59)? mem[548] : 
                         (N61)? mem[612] : 
                         (N63)? mem[676] : 
                         (N65)? mem[740] : 
                         (N67)? mem[804] : 
                         (N69)? mem[868] : 
                         (N71)? mem[932] : 
                         (N73)? mem[996] : 
                         (N44)? mem[1060] : 
                         (N46)? mem[1124] : 
                         (N48)? mem[1188] : 
                         (N50)? mem[1252] : 
                         (N52)? mem[1316] : 
                         (N54)? mem[1380] : 
                         (N56)? mem[1444] : 
                         (N58)? mem[1508] : 
                         (N60)? mem[1572] : 
                         (N62)? mem[1636] : 
                         (N64)? mem[1700] : 
                         (N66)? mem[1764] : 
                         (N68)? mem[1828] : 
                         (N70)? mem[1892] : 
                         (N72)? mem[1956] : 
                         (N74)? mem[2020] : 1'b0;
  assign r0_data_o[35] = (N43)? mem[35] : 
                         (N45)? mem[99] : 
                         (N47)? mem[163] : 
                         (N49)? mem[227] : 
                         (N51)? mem[291] : 
                         (N53)? mem[355] : 
                         (N55)? mem[419] : 
                         (N57)? mem[483] : 
                         (N59)? mem[547] : 
                         (N61)? mem[611] : 
                         (N63)? mem[675] : 
                         (N65)? mem[739] : 
                         (N67)? mem[803] : 
                         (N69)? mem[867] : 
                         (N71)? mem[931] : 
                         (N73)? mem[995] : 
                         (N44)? mem[1059] : 
                         (N46)? mem[1123] : 
                         (N48)? mem[1187] : 
                         (N50)? mem[1251] : 
                         (N52)? mem[1315] : 
                         (N54)? mem[1379] : 
                         (N56)? mem[1443] : 
                         (N58)? mem[1507] : 
                         (N60)? mem[1571] : 
                         (N62)? mem[1635] : 
                         (N64)? mem[1699] : 
                         (N66)? mem[1763] : 
                         (N68)? mem[1827] : 
                         (N70)? mem[1891] : 
                         (N72)? mem[1955] : 
                         (N74)? mem[2019] : 1'b0;
  assign r0_data_o[34] = (N43)? mem[34] : 
                         (N45)? mem[98] : 
                         (N47)? mem[162] : 
                         (N49)? mem[226] : 
                         (N51)? mem[290] : 
                         (N53)? mem[354] : 
                         (N55)? mem[418] : 
                         (N57)? mem[482] : 
                         (N59)? mem[546] : 
                         (N61)? mem[610] : 
                         (N63)? mem[674] : 
                         (N65)? mem[738] : 
                         (N67)? mem[802] : 
                         (N69)? mem[866] : 
                         (N71)? mem[930] : 
                         (N73)? mem[994] : 
                         (N44)? mem[1058] : 
                         (N46)? mem[1122] : 
                         (N48)? mem[1186] : 
                         (N50)? mem[1250] : 
                         (N52)? mem[1314] : 
                         (N54)? mem[1378] : 
                         (N56)? mem[1442] : 
                         (N58)? mem[1506] : 
                         (N60)? mem[1570] : 
                         (N62)? mem[1634] : 
                         (N64)? mem[1698] : 
                         (N66)? mem[1762] : 
                         (N68)? mem[1826] : 
                         (N70)? mem[1890] : 
                         (N72)? mem[1954] : 
                         (N74)? mem[2018] : 1'b0;
  assign r0_data_o[33] = (N43)? mem[33] : 
                         (N45)? mem[97] : 
                         (N47)? mem[161] : 
                         (N49)? mem[225] : 
                         (N51)? mem[289] : 
                         (N53)? mem[353] : 
                         (N55)? mem[417] : 
                         (N57)? mem[481] : 
                         (N59)? mem[545] : 
                         (N61)? mem[609] : 
                         (N63)? mem[673] : 
                         (N65)? mem[737] : 
                         (N67)? mem[801] : 
                         (N69)? mem[865] : 
                         (N71)? mem[929] : 
                         (N73)? mem[993] : 
                         (N44)? mem[1057] : 
                         (N46)? mem[1121] : 
                         (N48)? mem[1185] : 
                         (N50)? mem[1249] : 
                         (N52)? mem[1313] : 
                         (N54)? mem[1377] : 
                         (N56)? mem[1441] : 
                         (N58)? mem[1505] : 
                         (N60)? mem[1569] : 
                         (N62)? mem[1633] : 
                         (N64)? mem[1697] : 
                         (N66)? mem[1761] : 
                         (N68)? mem[1825] : 
                         (N70)? mem[1889] : 
                         (N72)? mem[1953] : 
                         (N74)? mem[2017] : 1'b0;
  assign r0_data_o[32] = (N43)? mem[32] : 
                         (N45)? mem[96] : 
                         (N47)? mem[160] : 
                         (N49)? mem[224] : 
                         (N51)? mem[288] : 
                         (N53)? mem[352] : 
                         (N55)? mem[416] : 
                         (N57)? mem[480] : 
                         (N59)? mem[544] : 
                         (N61)? mem[608] : 
                         (N63)? mem[672] : 
                         (N65)? mem[736] : 
                         (N67)? mem[800] : 
                         (N69)? mem[864] : 
                         (N71)? mem[928] : 
                         (N73)? mem[992] : 
                         (N44)? mem[1056] : 
                         (N46)? mem[1120] : 
                         (N48)? mem[1184] : 
                         (N50)? mem[1248] : 
                         (N52)? mem[1312] : 
                         (N54)? mem[1376] : 
                         (N56)? mem[1440] : 
                         (N58)? mem[1504] : 
                         (N60)? mem[1568] : 
                         (N62)? mem[1632] : 
                         (N64)? mem[1696] : 
                         (N66)? mem[1760] : 
                         (N68)? mem[1824] : 
                         (N70)? mem[1888] : 
                         (N72)? mem[1952] : 
                         (N74)? mem[2016] : 1'b0;
  assign r0_data_o[31] = (N43)? mem[31] : 
                         (N45)? mem[95] : 
                         (N47)? mem[159] : 
                         (N49)? mem[223] : 
                         (N51)? mem[287] : 
                         (N53)? mem[351] : 
                         (N55)? mem[415] : 
                         (N57)? mem[479] : 
                         (N59)? mem[543] : 
                         (N61)? mem[607] : 
                         (N63)? mem[671] : 
                         (N65)? mem[735] : 
                         (N67)? mem[799] : 
                         (N69)? mem[863] : 
                         (N71)? mem[927] : 
                         (N73)? mem[991] : 
                         (N44)? mem[1055] : 
                         (N46)? mem[1119] : 
                         (N48)? mem[1183] : 
                         (N50)? mem[1247] : 
                         (N52)? mem[1311] : 
                         (N54)? mem[1375] : 
                         (N56)? mem[1439] : 
                         (N58)? mem[1503] : 
                         (N60)? mem[1567] : 
                         (N62)? mem[1631] : 
                         (N64)? mem[1695] : 
                         (N66)? mem[1759] : 
                         (N68)? mem[1823] : 
                         (N70)? mem[1887] : 
                         (N72)? mem[1951] : 
                         (N74)? mem[2015] : 1'b0;
  assign r0_data_o[30] = (N43)? mem[30] : 
                         (N45)? mem[94] : 
                         (N47)? mem[158] : 
                         (N49)? mem[222] : 
                         (N51)? mem[286] : 
                         (N53)? mem[350] : 
                         (N55)? mem[414] : 
                         (N57)? mem[478] : 
                         (N59)? mem[542] : 
                         (N61)? mem[606] : 
                         (N63)? mem[670] : 
                         (N65)? mem[734] : 
                         (N67)? mem[798] : 
                         (N69)? mem[862] : 
                         (N71)? mem[926] : 
                         (N73)? mem[990] : 
                         (N44)? mem[1054] : 
                         (N46)? mem[1118] : 
                         (N48)? mem[1182] : 
                         (N50)? mem[1246] : 
                         (N52)? mem[1310] : 
                         (N54)? mem[1374] : 
                         (N56)? mem[1438] : 
                         (N58)? mem[1502] : 
                         (N60)? mem[1566] : 
                         (N62)? mem[1630] : 
                         (N64)? mem[1694] : 
                         (N66)? mem[1758] : 
                         (N68)? mem[1822] : 
                         (N70)? mem[1886] : 
                         (N72)? mem[1950] : 
                         (N74)? mem[2014] : 1'b0;
  assign r0_data_o[29] = (N43)? mem[29] : 
                         (N45)? mem[93] : 
                         (N47)? mem[157] : 
                         (N49)? mem[221] : 
                         (N51)? mem[285] : 
                         (N53)? mem[349] : 
                         (N55)? mem[413] : 
                         (N57)? mem[477] : 
                         (N59)? mem[541] : 
                         (N61)? mem[605] : 
                         (N63)? mem[669] : 
                         (N65)? mem[733] : 
                         (N67)? mem[797] : 
                         (N69)? mem[861] : 
                         (N71)? mem[925] : 
                         (N73)? mem[989] : 
                         (N44)? mem[1053] : 
                         (N46)? mem[1117] : 
                         (N48)? mem[1181] : 
                         (N50)? mem[1245] : 
                         (N52)? mem[1309] : 
                         (N54)? mem[1373] : 
                         (N56)? mem[1437] : 
                         (N58)? mem[1501] : 
                         (N60)? mem[1565] : 
                         (N62)? mem[1629] : 
                         (N64)? mem[1693] : 
                         (N66)? mem[1757] : 
                         (N68)? mem[1821] : 
                         (N70)? mem[1885] : 
                         (N72)? mem[1949] : 
                         (N74)? mem[2013] : 1'b0;
  assign r0_data_o[28] = (N43)? mem[28] : 
                         (N45)? mem[92] : 
                         (N47)? mem[156] : 
                         (N49)? mem[220] : 
                         (N51)? mem[284] : 
                         (N53)? mem[348] : 
                         (N55)? mem[412] : 
                         (N57)? mem[476] : 
                         (N59)? mem[540] : 
                         (N61)? mem[604] : 
                         (N63)? mem[668] : 
                         (N65)? mem[732] : 
                         (N67)? mem[796] : 
                         (N69)? mem[860] : 
                         (N71)? mem[924] : 
                         (N73)? mem[988] : 
                         (N44)? mem[1052] : 
                         (N46)? mem[1116] : 
                         (N48)? mem[1180] : 
                         (N50)? mem[1244] : 
                         (N52)? mem[1308] : 
                         (N54)? mem[1372] : 
                         (N56)? mem[1436] : 
                         (N58)? mem[1500] : 
                         (N60)? mem[1564] : 
                         (N62)? mem[1628] : 
                         (N64)? mem[1692] : 
                         (N66)? mem[1756] : 
                         (N68)? mem[1820] : 
                         (N70)? mem[1884] : 
                         (N72)? mem[1948] : 
                         (N74)? mem[2012] : 1'b0;
  assign r0_data_o[27] = (N43)? mem[27] : 
                         (N45)? mem[91] : 
                         (N47)? mem[155] : 
                         (N49)? mem[219] : 
                         (N51)? mem[283] : 
                         (N53)? mem[347] : 
                         (N55)? mem[411] : 
                         (N57)? mem[475] : 
                         (N59)? mem[539] : 
                         (N61)? mem[603] : 
                         (N63)? mem[667] : 
                         (N65)? mem[731] : 
                         (N67)? mem[795] : 
                         (N69)? mem[859] : 
                         (N71)? mem[923] : 
                         (N73)? mem[987] : 
                         (N44)? mem[1051] : 
                         (N46)? mem[1115] : 
                         (N48)? mem[1179] : 
                         (N50)? mem[1243] : 
                         (N52)? mem[1307] : 
                         (N54)? mem[1371] : 
                         (N56)? mem[1435] : 
                         (N58)? mem[1499] : 
                         (N60)? mem[1563] : 
                         (N62)? mem[1627] : 
                         (N64)? mem[1691] : 
                         (N66)? mem[1755] : 
                         (N68)? mem[1819] : 
                         (N70)? mem[1883] : 
                         (N72)? mem[1947] : 
                         (N74)? mem[2011] : 1'b0;
  assign r0_data_o[26] = (N43)? mem[26] : 
                         (N45)? mem[90] : 
                         (N47)? mem[154] : 
                         (N49)? mem[218] : 
                         (N51)? mem[282] : 
                         (N53)? mem[346] : 
                         (N55)? mem[410] : 
                         (N57)? mem[474] : 
                         (N59)? mem[538] : 
                         (N61)? mem[602] : 
                         (N63)? mem[666] : 
                         (N65)? mem[730] : 
                         (N67)? mem[794] : 
                         (N69)? mem[858] : 
                         (N71)? mem[922] : 
                         (N73)? mem[986] : 
                         (N44)? mem[1050] : 
                         (N46)? mem[1114] : 
                         (N48)? mem[1178] : 
                         (N50)? mem[1242] : 
                         (N52)? mem[1306] : 
                         (N54)? mem[1370] : 
                         (N56)? mem[1434] : 
                         (N58)? mem[1498] : 
                         (N60)? mem[1562] : 
                         (N62)? mem[1626] : 
                         (N64)? mem[1690] : 
                         (N66)? mem[1754] : 
                         (N68)? mem[1818] : 
                         (N70)? mem[1882] : 
                         (N72)? mem[1946] : 
                         (N74)? mem[2010] : 1'b0;
  assign r0_data_o[25] = (N43)? mem[25] : 
                         (N45)? mem[89] : 
                         (N47)? mem[153] : 
                         (N49)? mem[217] : 
                         (N51)? mem[281] : 
                         (N53)? mem[345] : 
                         (N55)? mem[409] : 
                         (N57)? mem[473] : 
                         (N59)? mem[537] : 
                         (N61)? mem[601] : 
                         (N63)? mem[665] : 
                         (N65)? mem[729] : 
                         (N67)? mem[793] : 
                         (N69)? mem[857] : 
                         (N71)? mem[921] : 
                         (N73)? mem[985] : 
                         (N44)? mem[1049] : 
                         (N46)? mem[1113] : 
                         (N48)? mem[1177] : 
                         (N50)? mem[1241] : 
                         (N52)? mem[1305] : 
                         (N54)? mem[1369] : 
                         (N56)? mem[1433] : 
                         (N58)? mem[1497] : 
                         (N60)? mem[1561] : 
                         (N62)? mem[1625] : 
                         (N64)? mem[1689] : 
                         (N66)? mem[1753] : 
                         (N68)? mem[1817] : 
                         (N70)? mem[1881] : 
                         (N72)? mem[1945] : 
                         (N74)? mem[2009] : 1'b0;
  assign r0_data_o[24] = (N43)? mem[24] : 
                         (N45)? mem[88] : 
                         (N47)? mem[152] : 
                         (N49)? mem[216] : 
                         (N51)? mem[280] : 
                         (N53)? mem[344] : 
                         (N55)? mem[408] : 
                         (N57)? mem[472] : 
                         (N59)? mem[536] : 
                         (N61)? mem[600] : 
                         (N63)? mem[664] : 
                         (N65)? mem[728] : 
                         (N67)? mem[792] : 
                         (N69)? mem[856] : 
                         (N71)? mem[920] : 
                         (N73)? mem[984] : 
                         (N44)? mem[1048] : 
                         (N46)? mem[1112] : 
                         (N48)? mem[1176] : 
                         (N50)? mem[1240] : 
                         (N52)? mem[1304] : 
                         (N54)? mem[1368] : 
                         (N56)? mem[1432] : 
                         (N58)? mem[1496] : 
                         (N60)? mem[1560] : 
                         (N62)? mem[1624] : 
                         (N64)? mem[1688] : 
                         (N66)? mem[1752] : 
                         (N68)? mem[1816] : 
                         (N70)? mem[1880] : 
                         (N72)? mem[1944] : 
                         (N74)? mem[2008] : 1'b0;
  assign r0_data_o[23] = (N43)? mem[23] : 
                         (N45)? mem[87] : 
                         (N47)? mem[151] : 
                         (N49)? mem[215] : 
                         (N51)? mem[279] : 
                         (N53)? mem[343] : 
                         (N55)? mem[407] : 
                         (N57)? mem[471] : 
                         (N59)? mem[535] : 
                         (N61)? mem[599] : 
                         (N63)? mem[663] : 
                         (N65)? mem[727] : 
                         (N67)? mem[791] : 
                         (N69)? mem[855] : 
                         (N71)? mem[919] : 
                         (N73)? mem[983] : 
                         (N44)? mem[1047] : 
                         (N46)? mem[1111] : 
                         (N48)? mem[1175] : 
                         (N50)? mem[1239] : 
                         (N52)? mem[1303] : 
                         (N54)? mem[1367] : 
                         (N56)? mem[1431] : 
                         (N58)? mem[1495] : 
                         (N60)? mem[1559] : 
                         (N62)? mem[1623] : 
                         (N64)? mem[1687] : 
                         (N66)? mem[1751] : 
                         (N68)? mem[1815] : 
                         (N70)? mem[1879] : 
                         (N72)? mem[1943] : 
                         (N74)? mem[2007] : 1'b0;
  assign r0_data_o[22] = (N43)? mem[22] : 
                         (N45)? mem[86] : 
                         (N47)? mem[150] : 
                         (N49)? mem[214] : 
                         (N51)? mem[278] : 
                         (N53)? mem[342] : 
                         (N55)? mem[406] : 
                         (N57)? mem[470] : 
                         (N59)? mem[534] : 
                         (N61)? mem[598] : 
                         (N63)? mem[662] : 
                         (N65)? mem[726] : 
                         (N67)? mem[790] : 
                         (N69)? mem[854] : 
                         (N71)? mem[918] : 
                         (N73)? mem[982] : 
                         (N44)? mem[1046] : 
                         (N46)? mem[1110] : 
                         (N48)? mem[1174] : 
                         (N50)? mem[1238] : 
                         (N52)? mem[1302] : 
                         (N54)? mem[1366] : 
                         (N56)? mem[1430] : 
                         (N58)? mem[1494] : 
                         (N60)? mem[1558] : 
                         (N62)? mem[1622] : 
                         (N64)? mem[1686] : 
                         (N66)? mem[1750] : 
                         (N68)? mem[1814] : 
                         (N70)? mem[1878] : 
                         (N72)? mem[1942] : 
                         (N74)? mem[2006] : 1'b0;
  assign r0_data_o[21] = (N43)? mem[21] : 
                         (N45)? mem[85] : 
                         (N47)? mem[149] : 
                         (N49)? mem[213] : 
                         (N51)? mem[277] : 
                         (N53)? mem[341] : 
                         (N55)? mem[405] : 
                         (N57)? mem[469] : 
                         (N59)? mem[533] : 
                         (N61)? mem[597] : 
                         (N63)? mem[661] : 
                         (N65)? mem[725] : 
                         (N67)? mem[789] : 
                         (N69)? mem[853] : 
                         (N71)? mem[917] : 
                         (N73)? mem[981] : 
                         (N44)? mem[1045] : 
                         (N46)? mem[1109] : 
                         (N48)? mem[1173] : 
                         (N50)? mem[1237] : 
                         (N52)? mem[1301] : 
                         (N54)? mem[1365] : 
                         (N56)? mem[1429] : 
                         (N58)? mem[1493] : 
                         (N60)? mem[1557] : 
                         (N62)? mem[1621] : 
                         (N64)? mem[1685] : 
                         (N66)? mem[1749] : 
                         (N68)? mem[1813] : 
                         (N70)? mem[1877] : 
                         (N72)? mem[1941] : 
                         (N74)? mem[2005] : 1'b0;
  assign r0_data_o[20] = (N43)? mem[20] : 
                         (N45)? mem[84] : 
                         (N47)? mem[148] : 
                         (N49)? mem[212] : 
                         (N51)? mem[276] : 
                         (N53)? mem[340] : 
                         (N55)? mem[404] : 
                         (N57)? mem[468] : 
                         (N59)? mem[532] : 
                         (N61)? mem[596] : 
                         (N63)? mem[660] : 
                         (N65)? mem[724] : 
                         (N67)? mem[788] : 
                         (N69)? mem[852] : 
                         (N71)? mem[916] : 
                         (N73)? mem[980] : 
                         (N44)? mem[1044] : 
                         (N46)? mem[1108] : 
                         (N48)? mem[1172] : 
                         (N50)? mem[1236] : 
                         (N52)? mem[1300] : 
                         (N54)? mem[1364] : 
                         (N56)? mem[1428] : 
                         (N58)? mem[1492] : 
                         (N60)? mem[1556] : 
                         (N62)? mem[1620] : 
                         (N64)? mem[1684] : 
                         (N66)? mem[1748] : 
                         (N68)? mem[1812] : 
                         (N70)? mem[1876] : 
                         (N72)? mem[1940] : 
                         (N74)? mem[2004] : 1'b0;
  assign r0_data_o[19] = (N43)? mem[19] : 
                         (N45)? mem[83] : 
                         (N47)? mem[147] : 
                         (N49)? mem[211] : 
                         (N51)? mem[275] : 
                         (N53)? mem[339] : 
                         (N55)? mem[403] : 
                         (N57)? mem[467] : 
                         (N59)? mem[531] : 
                         (N61)? mem[595] : 
                         (N63)? mem[659] : 
                         (N65)? mem[723] : 
                         (N67)? mem[787] : 
                         (N69)? mem[851] : 
                         (N71)? mem[915] : 
                         (N73)? mem[979] : 
                         (N44)? mem[1043] : 
                         (N46)? mem[1107] : 
                         (N48)? mem[1171] : 
                         (N50)? mem[1235] : 
                         (N52)? mem[1299] : 
                         (N54)? mem[1363] : 
                         (N56)? mem[1427] : 
                         (N58)? mem[1491] : 
                         (N60)? mem[1555] : 
                         (N62)? mem[1619] : 
                         (N64)? mem[1683] : 
                         (N66)? mem[1747] : 
                         (N68)? mem[1811] : 
                         (N70)? mem[1875] : 
                         (N72)? mem[1939] : 
                         (N74)? mem[2003] : 1'b0;
  assign r0_data_o[18] = (N43)? mem[18] : 
                         (N45)? mem[82] : 
                         (N47)? mem[146] : 
                         (N49)? mem[210] : 
                         (N51)? mem[274] : 
                         (N53)? mem[338] : 
                         (N55)? mem[402] : 
                         (N57)? mem[466] : 
                         (N59)? mem[530] : 
                         (N61)? mem[594] : 
                         (N63)? mem[658] : 
                         (N65)? mem[722] : 
                         (N67)? mem[786] : 
                         (N69)? mem[850] : 
                         (N71)? mem[914] : 
                         (N73)? mem[978] : 
                         (N44)? mem[1042] : 
                         (N46)? mem[1106] : 
                         (N48)? mem[1170] : 
                         (N50)? mem[1234] : 
                         (N52)? mem[1298] : 
                         (N54)? mem[1362] : 
                         (N56)? mem[1426] : 
                         (N58)? mem[1490] : 
                         (N60)? mem[1554] : 
                         (N62)? mem[1618] : 
                         (N64)? mem[1682] : 
                         (N66)? mem[1746] : 
                         (N68)? mem[1810] : 
                         (N70)? mem[1874] : 
                         (N72)? mem[1938] : 
                         (N74)? mem[2002] : 1'b0;
  assign r0_data_o[17] = (N43)? mem[17] : 
                         (N45)? mem[81] : 
                         (N47)? mem[145] : 
                         (N49)? mem[209] : 
                         (N51)? mem[273] : 
                         (N53)? mem[337] : 
                         (N55)? mem[401] : 
                         (N57)? mem[465] : 
                         (N59)? mem[529] : 
                         (N61)? mem[593] : 
                         (N63)? mem[657] : 
                         (N65)? mem[721] : 
                         (N67)? mem[785] : 
                         (N69)? mem[849] : 
                         (N71)? mem[913] : 
                         (N73)? mem[977] : 
                         (N44)? mem[1041] : 
                         (N46)? mem[1105] : 
                         (N48)? mem[1169] : 
                         (N50)? mem[1233] : 
                         (N52)? mem[1297] : 
                         (N54)? mem[1361] : 
                         (N56)? mem[1425] : 
                         (N58)? mem[1489] : 
                         (N60)? mem[1553] : 
                         (N62)? mem[1617] : 
                         (N64)? mem[1681] : 
                         (N66)? mem[1745] : 
                         (N68)? mem[1809] : 
                         (N70)? mem[1873] : 
                         (N72)? mem[1937] : 
                         (N74)? mem[2001] : 1'b0;
  assign r0_data_o[16] = (N43)? mem[16] : 
                         (N45)? mem[80] : 
                         (N47)? mem[144] : 
                         (N49)? mem[208] : 
                         (N51)? mem[272] : 
                         (N53)? mem[336] : 
                         (N55)? mem[400] : 
                         (N57)? mem[464] : 
                         (N59)? mem[528] : 
                         (N61)? mem[592] : 
                         (N63)? mem[656] : 
                         (N65)? mem[720] : 
                         (N67)? mem[784] : 
                         (N69)? mem[848] : 
                         (N71)? mem[912] : 
                         (N73)? mem[976] : 
                         (N44)? mem[1040] : 
                         (N46)? mem[1104] : 
                         (N48)? mem[1168] : 
                         (N50)? mem[1232] : 
                         (N52)? mem[1296] : 
                         (N54)? mem[1360] : 
                         (N56)? mem[1424] : 
                         (N58)? mem[1488] : 
                         (N60)? mem[1552] : 
                         (N62)? mem[1616] : 
                         (N64)? mem[1680] : 
                         (N66)? mem[1744] : 
                         (N68)? mem[1808] : 
                         (N70)? mem[1872] : 
                         (N72)? mem[1936] : 
                         (N74)? mem[2000] : 1'b0;
  assign r0_data_o[15] = (N43)? mem[15] : 
                         (N45)? mem[79] : 
                         (N47)? mem[143] : 
                         (N49)? mem[207] : 
                         (N51)? mem[271] : 
                         (N53)? mem[335] : 
                         (N55)? mem[399] : 
                         (N57)? mem[463] : 
                         (N59)? mem[527] : 
                         (N61)? mem[591] : 
                         (N63)? mem[655] : 
                         (N65)? mem[719] : 
                         (N67)? mem[783] : 
                         (N69)? mem[847] : 
                         (N71)? mem[911] : 
                         (N73)? mem[975] : 
                         (N44)? mem[1039] : 
                         (N46)? mem[1103] : 
                         (N48)? mem[1167] : 
                         (N50)? mem[1231] : 
                         (N52)? mem[1295] : 
                         (N54)? mem[1359] : 
                         (N56)? mem[1423] : 
                         (N58)? mem[1487] : 
                         (N60)? mem[1551] : 
                         (N62)? mem[1615] : 
                         (N64)? mem[1679] : 
                         (N66)? mem[1743] : 
                         (N68)? mem[1807] : 
                         (N70)? mem[1871] : 
                         (N72)? mem[1935] : 
                         (N74)? mem[1999] : 1'b0;
  assign r0_data_o[14] = (N43)? mem[14] : 
                         (N45)? mem[78] : 
                         (N47)? mem[142] : 
                         (N49)? mem[206] : 
                         (N51)? mem[270] : 
                         (N53)? mem[334] : 
                         (N55)? mem[398] : 
                         (N57)? mem[462] : 
                         (N59)? mem[526] : 
                         (N61)? mem[590] : 
                         (N63)? mem[654] : 
                         (N65)? mem[718] : 
                         (N67)? mem[782] : 
                         (N69)? mem[846] : 
                         (N71)? mem[910] : 
                         (N73)? mem[974] : 
                         (N44)? mem[1038] : 
                         (N46)? mem[1102] : 
                         (N48)? mem[1166] : 
                         (N50)? mem[1230] : 
                         (N52)? mem[1294] : 
                         (N54)? mem[1358] : 
                         (N56)? mem[1422] : 
                         (N58)? mem[1486] : 
                         (N60)? mem[1550] : 
                         (N62)? mem[1614] : 
                         (N64)? mem[1678] : 
                         (N66)? mem[1742] : 
                         (N68)? mem[1806] : 
                         (N70)? mem[1870] : 
                         (N72)? mem[1934] : 
                         (N74)? mem[1998] : 1'b0;
  assign r0_data_o[13] = (N43)? mem[13] : 
                         (N45)? mem[77] : 
                         (N47)? mem[141] : 
                         (N49)? mem[205] : 
                         (N51)? mem[269] : 
                         (N53)? mem[333] : 
                         (N55)? mem[397] : 
                         (N57)? mem[461] : 
                         (N59)? mem[525] : 
                         (N61)? mem[589] : 
                         (N63)? mem[653] : 
                         (N65)? mem[717] : 
                         (N67)? mem[781] : 
                         (N69)? mem[845] : 
                         (N71)? mem[909] : 
                         (N73)? mem[973] : 
                         (N44)? mem[1037] : 
                         (N46)? mem[1101] : 
                         (N48)? mem[1165] : 
                         (N50)? mem[1229] : 
                         (N52)? mem[1293] : 
                         (N54)? mem[1357] : 
                         (N56)? mem[1421] : 
                         (N58)? mem[1485] : 
                         (N60)? mem[1549] : 
                         (N62)? mem[1613] : 
                         (N64)? mem[1677] : 
                         (N66)? mem[1741] : 
                         (N68)? mem[1805] : 
                         (N70)? mem[1869] : 
                         (N72)? mem[1933] : 
                         (N74)? mem[1997] : 1'b0;
  assign r0_data_o[12] = (N43)? mem[12] : 
                         (N45)? mem[76] : 
                         (N47)? mem[140] : 
                         (N49)? mem[204] : 
                         (N51)? mem[268] : 
                         (N53)? mem[332] : 
                         (N55)? mem[396] : 
                         (N57)? mem[460] : 
                         (N59)? mem[524] : 
                         (N61)? mem[588] : 
                         (N63)? mem[652] : 
                         (N65)? mem[716] : 
                         (N67)? mem[780] : 
                         (N69)? mem[844] : 
                         (N71)? mem[908] : 
                         (N73)? mem[972] : 
                         (N44)? mem[1036] : 
                         (N46)? mem[1100] : 
                         (N48)? mem[1164] : 
                         (N50)? mem[1228] : 
                         (N52)? mem[1292] : 
                         (N54)? mem[1356] : 
                         (N56)? mem[1420] : 
                         (N58)? mem[1484] : 
                         (N60)? mem[1548] : 
                         (N62)? mem[1612] : 
                         (N64)? mem[1676] : 
                         (N66)? mem[1740] : 
                         (N68)? mem[1804] : 
                         (N70)? mem[1868] : 
                         (N72)? mem[1932] : 
                         (N74)? mem[1996] : 1'b0;
  assign r0_data_o[11] = (N43)? mem[11] : 
                         (N45)? mem[75] : 
                         (N47)? mem[139] : 
                         (N49)? mem[203] : 
                         (N51)? mem[267] : 
                         (N53)? mem[331] : 
                         (N55)? mem[395] : 
                         (N57)? mem[459] : 
                         (N59)? mem[523] : 
                         (N61)? mem[587] : 
                         (N63)? mem[651] : 
                         (N65)? mem[715] : 
                         (N67)? mem[779] : 
                         (N69)? mem[843] : 
                         (N71)? mem[907] : 
                         (N73)? mem[971] : 
                         (N44)? mem[1035] : 
                         (N46)? mem[1099] : 
                         (N48)? mem[1163] : 
                         (N50)? mem[1227] : 
                         (N52)? mem[1291] : 
                         (N54)? mem[1355] : 
                         (N56)? mem[1419] : 
                         (N58)? mem[1483] : 
                         (N60)? mem[1547] : 
                         (N62)? mem[1611] : 
                         (N64)? mem[1675] : 
                         (N66)? mem[1739] : 
                         (N68)? mem[1803] : 
                         (N70)? mem[1867] : 
                         (N72)? mem[1931] : 
                         (N74)? mem[1995] : 1'b0;
  assign r0_data_o[10] = (N43)? mem[10] : 
                         (N45)? mem[74] : 
                         (N47)? mem[138] : 
                         (N49)? mem[202] : 
                         (N51)? mem[266] : 
                         (N53)? mem[330] : 
                         (N55)? mem[394] : 
                         (N57)? mem[458] : 
                         (N59)? mem[522] : 
                         (N61)? mem[586] : 
                         (N63)? mem[650] : 
                         (N65)? mem[714] : 
                         (N67)? mem[778] : 
                         (N69)? mem[842] : 
                         (N71)? mem[906] : 
                         (N73)? mem[970] : 
                         (N44)? mem[1034] : 
                         (N46)? mem[1098] : 
                         (N48)? mem[1162] : 
                         (N50)? mem[1226] : 
                         (N52)? mem[1290] : 
                         (N54)? mem[1354] : 
                         (N56)? mem[1418] : 
                         (N58)? mem[1482] : 
                         (N60)? mem[1546] : 
                         (N62)? mem[1610] : 
                         (N64)? mem[1674] : 
                         (N66)? mem[1738] : 
                         (N68)? mem[1802] : 
                         (N70)? mem[1866] : 
                         (N72)? mem[1930] : 
                         (N74)? mem[1994] : 1'b0;
  assign r0_data_o[9] = (N43)? mem[9] : 
                        (N45)? mem[73] : 
                        (N47)? mem[137] : 
                        (N49)? mem[201] : 
                        (N51)? mem[265] : 
                        (N53)? mem[329] : 
                        (N55)? mem[393] : 
                        (N57)? mem[457] : 
                        (N59)? mem[521] : 
                        (N61)? mem[585] : 
                        (N63)? mem[649] : 
                        (N65)? mem[713] : 
                        (N67)? mem[777] : 
                        (N69)? mem[841] : 
                        (N71)? mem[905] : 
                        (N73)? mem[969] : 
                        (N44)? mem[1033] : 
                        (N46)? mem[1097] : 
                        (N48)? mem[1161] : 
                        (N50)? mem[1225] : 
                        (N52)? mem[1289] : 
                        (N54)? mem[1353] : 
                        (N56)? mem[1417] : 
                        (N58)? mem[1481] : 
                        (N60)? mem[1545] : 
                        (N62)? mem[1609] : 
                        (N64)? mem[1673] : 
                        (N66)? mem[1737] : 
                        (N68)? mem[1801] : 
                        (N70)? mem[1865] : 
                        (N72)? mem[1929] : 
                        (N74)? mem[1993] : 1'b0;
  assign r0_data_o[8] = (N43)? mem[8] : 
                        (N45)? mem[72] : 
                        (N47)? mem[136] : 
                        (N49)? mem[200] : 
                        (N51)? mem[264] : 
                        (N53)? mem[328] : 
                        (N55)? mem[392] : 
                        (N57)? mem[456] : 
                        (N59)? mem[520] : 
                        (N61)? mem[584] : 
                        (N63)? mem[648] : 
                        (N65)? mem[712] : 
                        (N67)? mem[776] : 
                        (N69)? mem[840] : 
                        (N71)? mem[904] : 
                        (N73)? mem[968] : 
                        (N44)? mem[1032] : 
                        (N46)? mem[1096] : 
                        (N48)? mem[1160] : 
                        (N50)? mem[1224] : 
                        (N52)? mem[1288] : 
                        (N54)? mem[1352] : 
                        (N56)? mem[1416] : 
                        (N58)? mem[1480] : 
                        (N60)? mem[1544] : 
                        (N62)? mem[1608] : 
                        (N64)? mem[1672] : 
                        (N66)? mem[1736] : 
                        (N68)? mem[1800] : 
                        (N70)? mem[1864] : 
                        (N72)? mem[1928] : 
                        (N74)? mem[1992] : 1'b0;
  assign r0_data_o[7] = (N43)? mem[7] : 
                        (N45)? mem[71] : 
                        (N47)? mem[135] : 
                        (N49)? mem[199] : 
                        (N51)? mem[263] : 
                        (N53)? mem[327] : 
                        (N55)? mem[391] : 
                        (N57)? mem[455] : 
                        (N59)? mem[519] : 
                        (N61)? mem[583] : 
                        (N63)? mem[647] : 
                        (N65)? mem[711] : 
                        (N67)? mem[775] : 
                        (N69)? mem[839] : 
                        (N71)? mem[903] : 
                        (N73)? mem[967] : 
                        (N44)? mem[1031] : 
                        (N46)? mem[1095] : 
                        (N48)? mem[1159] : 
                        (N50)? mem[1223] : 
                        (N52)? mem[1287] : 
                        (N54)? mem[1351] : 
                        (N56)? mem[1415] : 
                        (N58)? mem[1479] : 
                        (N60)? mem[1543] : 
                        (N62)? mem[1607] : 
                        (N64)? mem[1671] : 
                        (N66)? mem[1735] : 
                        (N68)? mem[1799] : 
                        (N70)? mem[1863] : 
                        (N72)? mem[1927] : 
                        (N74)? mem[1991] : 1'b0;
  assign r0_data_o[6] = (N43)? mem[6] : 
                        (N45)? mem[70] : 
                        (N47)? mem[134] : 
                        (N49)? mem[198] : 
                        (N51)? mem[262] : 
                        (N53)? mem[326] : 
                        (N55)? mem[390] : 
                        (N57)? mem[454] : 
                        (N59)? mem[518] : 
                        (N61)? mem[582] : 
                        (N63)? mem[646] : 
                        (N65)? mem[710] : 
                        (N67)? mem[774] : 
                        (N69)? mem[838] : 
                        (N71)? mem[902] : 
                        (N73)? mem[966] : 
                        (N44)? mem[1030] : 
                        (N46)? mem[1094] : 
                        (N48)? mem[1158] : 
                        (N50)? mem[1222] : 
                        (N52)? mem[1286] : 
                        (N54)? mem[1350] : 
                        (N56)? mem[1414] : 
                        (N58)? mem[1478] : 
                        (N60)? mem[1542] : 
                        (N62)? mem[1606] : 
                        (N64)? mem[1670] : 
                        (N66)? mem[1734] : 
                        (N68)? mem[1798] : 
                        (N70)? mem[1862] : 
                        (N72)? mem[1926] : 
                        (N74)? mem[1990] : 1'b0;
  assign r0_data_o[5] = (N43)? mem[5] : 
                        (N45)? mem[69] : 
                        (N47)? mem[133] : 
                        (N49)? mem[197] : 
                        (N51)? mem[261] : 
                        (N53)? mem[325] : 
                        (N55)? mem[389] : 
                        (N57)? mem[453] : 
                        (N59)? mem[517] : 
                        (N61)? mem[581] : 
                        (N63)? mem[645] : 
                        (N65)? mem[709] : 
                        (N67)? mem[773] : 
                        (N69)? mem[837] : 
                        (N71)? mem[901] : 
                        (N73)? mem[965] : 
                        (N44)? mem[1029] : 
                        (N46)? mem[1093] : 
                        (N48)? mem[1157] : 
                        (N50)? mem[1221] : 
                        (N52)? mem[1285] : 
                        (N54)? mem[1349] : 
                        (N56)? mem[1413] : 
                        (N58)? mem[1477] : 
                        (N60)? mem[1541] : 
                        (N62)? mem[1605] : 
                        (N64)? mem[1669] : 
                        (N66)? mem[1733] : 
                        (N68)? mem[1797] : 
                        (N70)? mem[1861] : 
                        (N72)? mem[1925] : 
                        (N74)? mem[1989] : 1'b0;
  assign r0_data_o[4] = (N43)? mem[4] : 
                        (N45)? mem[68] : 
                        (N47)? mem[132] : 
                        (N49)? mem[196] : 
                        (N51)? mem[260] : 
                        (N53)? mem[324] : 
                        (N55)? mem[388] : 
                        (N57)? mem[452] : 
                        (N59)? mem[516] : 
                        (N61)? mem[580] : 
                        (N63)? mem[644] : 
                        (N65)? mem[708] : 
                        (N67)? mem[772] : 
                        (N69)? mem[836] : 
                        (N71)? mem[900] : 
                        (N73)? mem[964] : 
                        (N44)? mem[1028] : 
                        (N46)? mem[1092] : 
                        (N48)? mem[1156] : 
                        (N50)? mem[1220] : 
                        (N52)? mem[1284] : 
                        (N54)? mem[1348] : 
                        (N56)? mem[1412] : 
                        (N58)? mem[1476] : 
                        (N60)? mem[1540] : 
                        (N62)? mem[1604] : 
                        (N64)? mem[1668] : 
                        (N66)? mem[1732] : 
                        (N68)? mem[1796] : 
                        (N70)? mem[1860] : 
                        (N72)? mem[1924] : 
                        (N74)? mem[1988] : 1'b0;
  assign r0_data_o[3] = (N43)? mem[3] : 
                        (N45)? mem[67] : 
                        (N47)? mem[131] : 
                        (N49)? mem[195] : 
                        (N51)? mem[259] : 
                        (N53)? mem[323] : 
                        (N55)? mem[387] : 
                        (N57)? mem[451] : 
                        (N59)? mem[515] : 
                        (N61)? mem[579] : 
                        (N63)? mem[643] : 
                        (N65)? mem[707] : 
                        (N67)? mem[771] : 
                        (N69)? mem[835] : 
                        (N71)? mem[899] : 
                        (N73)? mem[963] : 
                        (N44)? mem[1027] : 
                        (N46)? mem[1091] : 
                        (N48)? mem[1155] : 
                        (N50)? mem[1219] : 
                        (N52)? mem[1283] : 
                        (N54)? mem[1347] : 
                        (N56)? mem[1411] : 
                        (N58)? mem[1475] : 
                        (N60)? mem[1539] : 
                        (N62)? mem[1603] : 
                        (N64)? mem[1667] : 
                        (N66)? mem[1731] : 
                        (N68)? mem[1795] : 
                        (N70)? mem[1859] : 
                        (N72)? mem[1923] : 
                        (N74)? mem[1987] : 1'b0;
  assign r0_data_o[2] = (N43)? mem[2] : 
                        (N45)? mem[66] : 
                        (N47)? mem[130] : 
                        (N49)? mem[194] : 
                        (N51)? mem[258] : 
                        (N53)? mem[322] : 
                        (N55)? mem[386] : 
                        (N57)? mem[450] : 
                        (N59)? mem[514] : 
                        (N61)? mem[578] : 
                        (N63)? mem[642] : 
                        (N65)? mem[706] : 
                        (N67)? mem[770] : 
                        (N69)? mem[834] : 
                        (N71)? mem[898] : 
                        (N73)? mem[962] : 
                        (N44)? mem[1026] : 
                        (N46)? mem[1090] : 
                        (N48)? mem[1154] : 
                        (N50)? mem[1218] : 
                        (N52)? mem[1282] : 
                        (N54)? mem[1346] : 
                        (N56)? mem[1410] : 
                        (N58)? mem[1474] : 
                        (N60)? mem[1538] : 
                        (N62)? mem[1602] : 
                        (N64)? mem[1666] : 
                        (N66)? mem[1730] : 
                        (N68)? mem[1794] : 
                        (N70)? mem[1858] : 
                        (N72)? mem[1922] : 
                        (N74)? mem[1986] : 1'b0;
  assign r0_data_o[1] = (N43)? mem[1] : 
                        (N45)? mem[65] : 
                        (N47)? mem[129] : 
                        (N49)? mem[193] : 
                        (N51)? mem[257] : 
                        (N53)? mem[321] : 
                        (N55)? mem[385] : 
                        (N57)? mem[449] : 
                        (N59)? mem[513] : 
                        (N61)? mem[577] : 
                        (N63)? mem[641] : 
                        (N65)? mem[705] : 
                        (N67)? mem[769] : 
                        (N69)? mem[833] : 
                        (N71)? mem[897] : 
                        (N73)? mem[961] : 
                        (N44)? mem[1025] : 
                        (N46)? mem[1089] : 
                        (N48)? mem[1153] : 
                        (N50)? mem[1217] : 
                        (N52)? mem[1281] : 
                        (N54)? mem[1345] : 
                        (N56)? mem[1409] : 
                        (N58)? mem[1473] : 
                        (N60)? mem[1537] : 
                        (N62)? mem[1601] : 
                        (N64)? mem[1665] : 
                        (N66)? mem[1729] : 
                        (N68)? mem[1793] : 
                        (N70)? mem[1857] : 
                        (N72)? mem[1921] : 
                        (N74)? mem[1985] : 1'b0;
  assign r0_data_o[0] = (N43)? mem[0] : 
                        (N45)? mem[64] : 
                        (N47)? mem[128] : 
                        (N49)? mem[192] : 
                        (N51)? mem[256] : 
                        (N53)? mem[320] : 
                        (N55)? mem[384] : 
                        (N57)? mem[448] : 
                        (N59)? mem[512] : 
                        (N61)? mem[576] : 
                        (N63)? mem[640] : 
                        (N65)? mem[704] : 
                        (N67)? mem[768] : 
                        (N69)? mem[832] : 
                        (N71)? mem[896] : 
                        (N73)? mem[960] : 
                        (N44)? mem[1024] : 
                        (N46)? mem[1088] : 
                        (N48)? mem[1152] : 
                        (N50)? mem[1216] : 
                        (N52)? mem[1280] : 
                        (N54)? mem[1344] : 
                        (N56)? mem[1408] : 
                        (N58)? mem[1472] : 
                        (N60)? mem[1536] : 
                        (N62)? mem[1600] : 
                        (N64)? mem[1664] : 
                        (N66)? mem[1728] : 
                        (N68)? mem[1792] : 
                        (N70)? mem[1856] : 
                        (N72)? mem[1920] : 
                        (N74)? mem[1984] : 1'b0;
  assign r1_data_o[63] = (N108)? mem[63] : 
                         (N110)? mem[127] : 
                         (N112)? mem[191] : 
                         (N114)? mem[255] : 
                         (N116)? mem[319] : 
                         (N118)? mem[383] : 
                         (N120)? mem[447] : 
                         (N122)? mem[511] : 
                         (N124)? mem[575] : 
                         (N126)? mem[639] : 
                         (N128)? mem[703] : 
                         (N130)? mem[767] : 
                         (N132)? mem[831] : 
                         (N134)? mem[895] : 
                         (N136)? mem[959] : 
                         (N138)? mem[1023] : 
                         (N109)? mem[1087] : 
                         (N111)? mem[1151] : 
                         (N113)? mem[1215] : 
                         (N115)? mem[1279] : 
                         (N117)? mem[1343] : 
                         (N119)? mem[1407] : 
                         (N121)? mem[1471] : 
                         (N123)? mem[1535] : 
                         (N125)? mem[1599] : 
                         (N127)? mem[1663] : 
                         (N129)? mem[1727] : 
                         (N131)? mem[1791] : 
                         (N133)? mem[1855] : 
                         (N135)? mem[1919] : 
                         (N137)? mem[1983] : 
                         (N139)? mem[2047] : 1'b0;
  assign r1_data_o[62] = (N108)? mem[62] : 
                         (N110)? mem[126] : 
                         (N112)? mem[190] : 
                         (N114)? mem[254] : 
                         (N116)? mem[318] : 
                         (N118)? mem[382] : 
                         (N120)? mem[446] : 
                         (N122)? mem[510] : 
                         (N124)? mem[574] : 
                         (N126)? mem[638] : 
                         (N128)? mem[702] : 
                         (N130)? mem[766] : 
                         (N132)? mem[830] : 
                         (N134)? mem[894] : 
                         (N136)? mem[958] : 
                         (N138)? mem[1022] : 
                         (N109)? mem[1086] : 
                         (N111)? mem[1150] : 
                         (N113)? mem[1214] : 
                         (N115)? mem[1278] : 
                         (N117)? mem[1342] : 
                         (N119)? mem[1406] : 
                         (N121)? mem[1470] : 
                         (N123)? mem[1534] : 
                         (N125)? mem[1598] : 
                         (N127)? mem[1662] : 
                         (N129)? mem[1726] : 
                         (N131)? mem[1790] : 
                         (N133)? mem[1854] : 
                         (N135)? mem[1918] : 
                         (N137)? mem[1982] : 
                         (N139)? mem[2046] : 1'b0;
  assign r1_data_o[61] = (N108)? mem[61] : 
                         (N110)? mem[125] : 
                         (N112)? mem[189] : 
                         (N114)? mem[253] : 
                         (N116)? mem[317] : 
                         (N118)? mem[381] : 
                         (N120)? mem[445] : 
                         (N122)? mem[509] : 
                         (N124)? mem[573] : 
                         (N126)? mem[637] : 
                         (N128)? mem[701] : 
                         (N130)? mem[765] : 
                         (N132)? mem[829] : 
                         (N134)? mem[893] : 
                         (N136)? mem[957] : 
                         (N138)? mem[1021] : 
                         (N109)? mem[1085] : 
                         (N111)? mem[1149] : 
                         (N113)? mem[1213] : 
                         (N115)? mem[1277] : 
                         (N117)? mem[1341] : 
                         (N119)? mem[1405] : 
                         (N121)? mem[1469] : 
                         (N123)? mem[1533] : 
                         (N125)? mem[1597] : 
                         (N127)? mem[1661] : 
                         (N129)? mem[1725] : 
                         (N131)? mem[1789] : 
                         (N133)? mem[1853] : 
                         (N135)? mem[1917] : 
                         (N137)? mem[1981] : 
                         (N139)? mem[2045] : 1'b0;
  assign r1_data_o[60] = (N108)? mem[60] : 
                         (N110)? mem[124] : 
                         (N112)? mem[188] : 
                         (N114)? mem[252] : 
                         (N116)? mem[316] : 
                         (N118)? mem[380] : 
                         (N120)? mem[444] : 
                         (N122)? mem[508] : 
                         (N124)? mem[572] : 
                         (N126)? mem[636] : 
                         (N128)? mem[700] : 
                         (N130)? mem[764] : 
                         (N132)? mem[828] : 
                         (N134)? mem[892] : 
                         (N136)? mem[956] : 
                         (N138)? mem[1020] : 
                         (N109)? mem[1084] : 
                         (N111)? mem[1148] : 
                         (N113)? mem[1212] : 
                         (N115)? mem[1276] : 
                         (N117)? mem[1340] : 
                         (N119)? mem[1404] : 
                         (N121)? mem[1468] : 
                         (N123)? mem[1532] : 
                         (N125)? mem[1596] : 
                         (N127)? mem[1660] : 
                         (N129)? mem[1724] : 
                         (N131)? mem[1788] : 
                         (N133)? mem[1852] : 
                         (N135)? mem[1916] : 
                         (N137)? mem[1980] : 
                         (N139)? mem[2044] : 1'b0;
  assign r1_data_o[59] = (N108)? mem[59] : 
                         (N110)? mem[123] : 
                         (N112)? mem[187] : 
                         (N114)? mem[251] : 
                         (N116)? mem[315] : 
                         (N118)? mem[379] : 
                         (N120)? mem[443] : 
                         (N122)? mem[507] : 
                         (N124)? mem[571] : 
                         (N126)? mem[635] : 
                         (N128)? mem[699] : 
                         (N130)? mem[763] : 
                         (N132)? mem[827] : 
                         (N134)? mem[891] : 
                         (N136)? mem[955] : 
                         (N138)? mem[1019] : 
                         (N109)? mem[1083] : 
                         (N111)? mem[1147] : 
                         (N113)? mem[1211] : 
                         (N115)? mem[1275] : 
                         (N117)? mem[1339] : 
                         (N119)? mem[1403] : 
                         (N121)? mem[1467] : 
                         (N123)? mem[1531] : 
                         (N125)? mem[1595] : 
                         (N127)? mem[1659] : 
                         (N129)? mem[1723] : 
                         (N131)? mem[1787] : 
                         (N133)? mem[1851] : 
                         (N135)? mem[1915] : 
                         (N137)? mem[1979] : 
                         (N139)? mem[2043] : 1'b0;
  assign r1_data_o[58] = (N108)? mem[58] : 
                         (N110)? mem[122] : 
                         (N112)? mem[186] : 
                         (N114)? mem[250] : 
                         (N116)? mem[314] : 
                         (N118)? mem[378] : 
                         (N120)? mem[442] : 
                         (N122)? mem[506] : 
                         (N124)? mem[570] : 
                         (N126)? mem[634] : 
                         (N128)? mem[698] : 
                         (N130)? mem[762] : 
                         (N132)? mem[826] : 
                         (N134)? mem[890] : 
                         (N136)? mem[954] : 
                         (N138)? mem[1018] : 
                         (N109)? mem[1082] : 
                         (N111)? mem[1146] : 
                         (N113)? mem[1210] : 
                         (N115)? mem[1274] : 
                         (N117)? mem[1338] : 
                         (N119)? mem[1402] : 
                         (N121)? mem[1466] : 
                         (N123)? mem[1530] : 
                         (N125)? mem[1594] : 
                         (N127)? mem[1658] : 
                         (N129)? mem[1722] : 
                         (N131)? mem[1786] : 
                         (N133)? mem[1850] : 
                         (N135)? mem[1914] : 
                         (N137)? mem[1978] : 
                         (N139)? mem[2042] : 1'b0;
  assign r1_data_o[57] = (N108)? mem[57] : 
                         (N110)? mem[121] : 
                         (N112)? mem[185] : 
                         (N114)? mem[249] : 
                         (N116)? mem[313] : 
                         (N118)? mem[377] : 
                         (N120)? mem[441] : 
                         (N122)? mem[505] : 
                         (N124)? mem[569] : 
                         (N126)? mem[633] : 
                         (N128)? mem[697] : 
                         (N130)? mem[761] : 
                         (N132)? mem[825] : 
                         (N134)? mem[889] : 
                         (N136)? mem[953] : 
                         (N138)? mem[1017] : 
                         (N109)? mem[1081] : 
                         (N111)? mem[1145] : 
                         (N113)? mem[1209] : 
                         (N115)? mem[1273] : 
                         (N117)? mem[1337] : 
                         (N119)? mem[1401] : 
                         (N121)? mem[1465] : 
                         (N123)? mem[1529] : 
                         (N125)? mem[1593] : 
                         (N127)? mem[1657] : 
                         (N129)? mem[1721] : 
                         (N131)? mem[1785] : 
                         (N133)? mem[1849] : 
                         (N135)? mem[1913] : 
                         (N137)? mem[1977] : 
                         (N139)? mem[2041] : 1'b0;
  assign r1_data_o[56] = (N108)? mem[56] : 
                         (N110)? mem[120] : 
                         (N112)? mem[184] : 
                         (N114)? mem[248] : 
                         (N116)? mem[312] : 
                         (N118)? mem[376] : 
                         (N120)? mem[440] : 
                         (N122)? mem[504] : 
                         (N124)? mem[568] : 
                         (N126)? mem[632] : 
                         (N128)? mem[696] : 
                         (N130)? mem[760] : 
                         (N132)? mem[824] : 
                         (N134)? mem[888] : 
                         (N136)? mem[952] : 
                         (N138)? mem[1016] : 
                         (N109)? mem[1080] : 
                         (N111)? mem[1144] : 
                         (N113)? mem[1208] : 
                         (N115)? mem[1272] : 
                         (N117)? mem[1336] : 
                         (N119)? mem[1400] : 
                         (N121)? mem[1464] : 
                         (N123)? mem[1528] : 
                         (N125)? mem[1592] : 
                         (N127)? mem[1656] : 
                         (N129)? mem[1720] : 
                         (N131)? mem[1784] : 
                         (N133)? mem[1848] : 
                         (N135)? mem[1912] : 
                         (N137)? mem[1976] : 
                         (N139)? mem[2040] : 1'b0;
  assign r1_data_o[55] = (N108)? mem[55] : 
                         (N110)? mem[119] : 
                         (N112)? mem[183] : 
                         (N114)? mem[247] : 
                         (N116)? mem[311] : 
                         (N118)? mem[375] : 
                         (N120)? mem[439] : 
                         (N122)? mem[503] : 
                         (N124)? mem[567] : 
                         (N126)? mem[631] : 
                         (N128)? mem[695] : 
                         (N130)? mem[759] : 
                         (N132)? mem[823] : 
                         (N134)? mem[887] : 
                         (N136)? mem[951] : 
                         (N138)? mem[1015] : 
                         (N109)? mem[1079] : 
                         (N111)? mem[1143] : 
                         (N113)? mem[1207] : 
                         (N115)? mem[1271] : 
                         (N117)? mem[1335] : 
                         (N119)? mem[1399] : 
                         (N121)? mem[1463] : 
                         (N123)? mem[1527] : 
                         (N125)? mem[1591] : 
                         (N127)? mem[1655] : 
                         (N129)? mem[1719] : 
                         (N131)? mem[1783] : 
                         (N133)? mem[1847] : 
                         (N135)? mem[1911] : 
                         (N137)? mem[1975] : 
                         (N139)? mem[2039] : 1'b0;
  assign r1_data_o[54] = (N108)? mem[54] : 
                         (N110)? mem[118] : 
                         (N112)? mem[182] : 
                         (N114)? mem[246] : 
                         (N116)? mem[310] : 
                         (N118)? mem[374] : 
                         (N120)? mem[438] : 
                         (N122)? mem[502] : 
                         (N124)? mem[566] : 
                         (N126)? mem[630] : 
                         (N128)? mem[694] : 
                         (N130)? mem[758] : 
                         (N132)? mem[822] : 
                         (N134)? mem[886] : 
                         (N136)? mem[950] : 
                         (N138)? mem[1014] : 
                         (N109)? mem[1078] : 
                         (N111)? mem[1142] : 
                         (N113)? mem[1206] : 
                         (N115)? mem[1270] : 
                         (N117)? mem[1334] : 
                         (N119)? mem[1398] : 
                         (N121)? mem[1462] : 
                         (N123)? mem[1526] : 
                         (N125)? mem[1590] : 
                         (N127)? mem[1654] : 
                         (N129)? mem[1718] : 
                         (N131)? mem[1782] : 
                         (N133)? mem[1846] : 
                         (N135)? mem[1910] : 
                         (N137)? mem[1974] : 
                         (N139)? mem[2038] : 1'b0;
  assign r1_data_o[53] = (N108)? mem[53] : 
                         (N110)? mem[117] : 
                         (N112)? mem[181] : 
                         (N114)? mem[245] : 
                         (N116)? mem[309] : 
                         (N118)? mem[373] : 
                         (N120)? mem[437] : 
                         (N122)? mem[501] : 
                         (N124)? mem[565] : 
                         (N126)? mem[629] : 
                         (N128)? mem[693] : 
                         (N130)? mem[757] : 
                         (N132)? mem[821] : 
                         (N134)? mem[885] : 
                         (N136)? mem[949] : 
                         (N138)? mem[1013] : 
                         (N109)? mem[1077] : 
                         (N111)? mem[1141] : 
                         (N113)? mem[1205] : 
                         (N115)? mem[1269] : 
                         (N117)? mem[1333] : 
                         (N119)? mem[1397] : 
                         (N121)? mem[1461] : 
                         (N123)? mem[1525] : 
                         (N125)? mem[1589] : 
                         (N127)? mem[1653] : 
                         (N129)? mem[1717] : 
                         (N131)? mem[1781] : 
                         (N133)? mem[1845] : 
                         (N135)? mem[1909] : 
                         (N137)? mem[1973] : 
                         (N139)? mem[2037] : 1'b0;
  assign r1_data_o[52] = (N108)? mem[52] : 
                         (N110)? mem[116] : 
                         (N112)? mem[180] : 
                         (N114)? mem[244] : 
                         (N116)? mem[308] : 
                         (N118)? mem[372] : 
                         (N120)? mem[436] : 
                         (N122)? mem[500] : 
                         (N124)? mem[564] : 
                         (N126)? mem[628] : 
                         (N128)? mem[692] : 
                         (N130)? mem[756] : 
                         (N132)? mem[820] : 
                         (N134)? mem[884] : 
                         (N136)? mem[948] : 
                         (N138)? mem[1012] : 
                         (N109)? mem[1076] : 
                         (N111)? mem[1140] : 
                         (N113)? mem[1204] : 
                         (N115)? mem[1268] : 
                         (N117)? mem[1332] : 
                         (N119)? mem[1396] : 
                         (N121)? mem[1460] : 
                         (N123)? mem[1524] : 
                         (N125)? mem[1588] : 
                         (N127)? mem[1652] : 
                         (N129)? mem[1716] : 
                         (N131)? mem[1780] : 
                         (N133)? mem[1844] : 
                         (N135)? mem[1908] : 
                         (N137)? mem[1972] : 
                         (N139)? mem[2036] : 1'b0;
  assign r1_data_o[51] = (N108)? mem[51] : 
                         (N110)? mem[115] : 
                         (N112)? mem[179] : 
                         (N114)? mem[243] : 
                         (N116)? mem[307] : 
                         (N118)? mem[371] : 
                         (N120)? mem[435] : 
                         (N122)? mem[499] : 
                         (N124)? mem[563] : 
                         (N126)? mem[627] : 
                         (N128)? mem[691] : 
                         (N130)? mem[755] : 
                         (N132)? mem[819] : 
                         (N134)? mem[883] : 
                         (N136)? mem[947] : 
                         (N138)? mem[1011] : 
                         (N109)? mem[1075] : 
                         (N111)? mem[1139] : 
                         (N113)? mem[1203] : 
                         (N115)? mem[1267] : 
                         (N117)? mem[1331] : 
                         (N119)? mem[1395] : 
                         (N121)? mem[1459] : 
                         (N123)? mem[1523] : 
                         (N125)? mem[1587] : 
                         (N127)? mem[1651] : 
                         (N129)? mem[1715] : 
                         (N131)? mem[1779] : 
                         (N133)? mem[1843] : 
                         (N135)? mem[1907] : 
                         (N137)? mem[1971] : 
                         (N139)? mem[2035] : 1'b0;
  assign r1_data_o[50] = (N108)? mem[50] : 
                         (N110)? mem[114] : 
                         (N112)? mem[178] : 
                         (N114)? mem[242] : 
                         (N116)? mem[306] : 
                         (N118)? mem[370] : 
                         (N120)? mem[434] : 
                         (N122)? mem[498] : 
                         (N124)? mem[562] : 
                         (N126)? mem[626] : 
                         (N128)? mem[690] : 
                         (N130)? mem[754] : 
                         (N132)? mem[818] : 
                         (N134)? mem[882] : 
                         (N136)? mem[946] : 
                         (N138)? mem[1010] : 
                         (N109)? mem[1074] : 
                         (N111)? mem[1138] : 
                         (N113)? mem[1202] : 
                         (N115)? mem[1266] : 
                         (N117)? mem[1330] : 
                         (N119)? mem[1394] : 
                         (N121)? mem[1458] : 
                         (N123)? mem[1522] : 
                         (N125)? mem[1586] : 
                         (N127)? mem[1650] : 
                         (N129)? mem[1714] : 
                         (N131)? mem[1778] : 
                         (N133)? mem[1842] : 
                         (N135)? mem[1906] : 
                         (N137)? mem[1970] : 
                         (N139)? mem[2034] : 1'b0;
  assign r1_data_o[49] = (N108)? mem[49] : 
                         (N110)? mem[113] : 
                         (N112)? mem[177] : 
                         (N114)? mem[241] : 
                         (N116)? mem[305] : 
                         (N118)? mem[369] : 
                         (N120)? mem[433] : 
                         (N122)? mem[497] : 
                         (N124)? mem[561] : 
                         (N126)? mem[625] : 
                         (N128)? mem[689] : 
                         (N130)? mem[753] : 
                         (N132)? mem[817] : 
                         (N134)? mem[881] : 
                         (N136)? mem[945] : 
                         (N138)? mem[1009] : 
                         (N109)? mem[1073] : 
                         (N111)? mem[1137] : 
                         (N113)? mem[1201] : 
                         (N115)? mem[1265] : 
                         (N117)? mem[1329] : 
                         (N119)? mem[1393] : 
                         (N121)? mem[1457] : 
                         (N123)? mem[1521] : 
                         (N125)? mem[1585] : 
                         (N127)? mem[1649] : 
                         (N129)? mem[1713] : 
                         (N131)? mem[1777] : 
                         (N133)? mem[1841] : 
                         (N135)? mem[1905] : 
                         (N137)? mem[1969] : 
                         (N139)? mem[2033] : 1'b0;
  assign r1_data_o[48] = (N108)? mem[48] : 
                         (N110)? mem[112] : 
                         (N112)? mem[176] : 
                         (N114)? mem[240] : 
                         (N116)? mem[304] : 
                         (N118)? mem[368] : 
                         (N120)? mem[432] : 
                         (N122)? mem[496] : 
                         (N124)? mem[560] : 
                         (N126)? mem[624] : 
                         (N128)? mem[688] : 
                         (N130)? mem[752] : 
                         (N132)? mem[816] : 
                         (N134)? mem[880] : 
                         (N136)? mem[944] : 
                         (N138)? mem[1008] : 
                         (N109)? mem[1072] : 
                         (N111)? mem[1136] : 
                         (N113)? mem[1200] : 
                         (N115)? mem[1264] : 
                         (N117)? mem[1328] : 
                         (N119)? mem[1392] : 
                         (N121)? mem[1456] : 
                         (N123)? mem[1520] : 
                         (N125)? mem[1584] : 
                         (N127)? mem[1648] : 
                         (N129)? mem[1712] : 
                         (N131)? mem[1776] : 
                         (N133)? mem[1840] : 
                         (N135)? mem[1904] : 
                         (N137)? mem[1968] : 
                         (N139)? mem[2032] : 1'b0;
  assign r1_data_o[47] = (N108)? mem[47] : 
                         (N110)? mem[111] : 
                         (N112)? mem[175] : 
                         (N114)? mem[239] : 
                         (N116)? mem[303] : 
                         (N118)? mem[367] : 
                         (N120)? mem[431] : 
                         (N122)? mem[495] : 
                         (N124)? mem[559] : 
                         (N126)? mem[623] : 
                         (N128)? mem[687] : 
                         (N130)? mem[751] : 
                         (N132)? mem[815] : 
                         (N134)? mem[879] : 
                         (N136)? mem[943] : 
                         (N138)? mem[1007] : 
                         (N109)? mem[1071] : 
                         (N111)? mem[1135] : 
                         (N113)? mem[1199] : 
                         (N115)? mem[1263] : 
                         (N117)? mem[1327] : 
                         (N119)? mem[1391] : 
                         (N121)? mem[1455] : 
                         (N123)? mem[1519] : 
                         (N125)? mem[1583] : 
                         (N127)? mem[1647] : 
                         (N129)? mem[1711] : 
                         (N131)? mem[1775] : 
                         (N133)? mem[1839] : 
                         (N135)? mem[1903] : 
                         (N137)? mem[1967] : 
                         (N139)? mem[2031] : 1'b0;
  assign r1_data_o[46] = (N108)? mem[46] : 
                         (N110)? mem[110] : 
                         (N112)? mem[174] : 
                         (N114)? mem[238] : 
                         (N116)? mem[302] : 
                         (N118)? mem[366] : 
                         (N120)? mem[430] : 
                         (N122)? mem[494] : 
                         (N124)? mem[558] : 
                         (N126)? mem[622] : 
                         (N128)? mem[686] : 
                         (N130)? mem[750] : 
                         (N132)? mem[814] : 
                         (N134)? mem[878] : 
                         (N136)? mem[942] : 
                         (N138)? mem[1006] : 
                         (N109)? mem[1070] : 
                         (N111)? mem[1134] : 
                         (N113)? mem[1198] : 
                         (N115)? mem[1262] : 
                         (N117)? mem[1326] : 
                         (N119)? mem[1390] : 
                         (N121)? mem[1454] : 
                         (N123)? mem[1518] : 
                         (N125)? mem[1582] : 
                         (N127)? mem[1646] : 
                         (N129)? mem[1710] : 
                         (N131)? mem[1774] : 
                         (N133)? mem[1838] : 
                         (N135)? mem[1902] : 
                         (N137)? mem[1966] : 
                         (N139)? mem[2030] : 1'b0;
  assign r1_data_o[45] = (N108)? mem[45] : 
                         (N110)? mem[109] : 
                         (N112)? mem[173] : 
                         (N114)? mem[237] : 
                         (N116)? mem[301] : 
                         (N118)? mem[365] : 
                         (N120)? mem[429] : 
                         (N122)? mem[493] : 
                         (N124)? mem[557] : 
                         (N126)? mem[621] : 
                         (N128)? mem[685] : 
                         (N130)? mem[749] : 
                         (N132)? mem[813] : 
                         (N134)? mem[877] : 
                         (N136)? mem[941] : 
                         (N138)? mem[1005] : 
                         (N109)? mem[1069] : 
                         (N111)? mem[1133] : 
                         (N113)? mem[1197] : 
                         (N115)? mem[1261] : 
                         (N117)? mem[1325] : 
                         (N119)? mem[1389] : 
                         (N121)? mem[1453] : 
                         (N123)? mem[1517] : 
                         (N125)? mem[1581] : 
                         (N127)? mem[1645] : 
                         (N129)? mem[1709] : 
                         (N131)? mem[1773] : 
                         (N133)? mem[1837] : 
                         (N135)? mem[1901] : 
                         (N137)? mem[1965] : 
                         (N139)? mem[2029] : 1'b0;
  assign r1_data_o[44] = (N108)? mem[44] : 
                         (N110)? mem[108] : 
                         (N112)? mem[172] : 
                         (N114)? mem[236] : 
                         (N116)? mem[300] : 
                         (N118)? mem[364] : 
                         (N120)? mem[428] : 
                         (N122)? mem[492] : 
                         (N124)? mem[556] : 
                         (N126)? mem[620] : 
                         (N128)? mem[684] : 
                         (N130)? mem[748] : 
                         (N132)? mem[812] : 
                         (N134)? mem[876] : 
                         (N136)? mem[940] : 
                         (N138)? mem[1004] : 
                         (N109)? mem[1068] : 
                         (N111)? mem[1132] : 
                         (N113)? mem[1196] : 
                         (N115)? mem[1260] : 
                         (N117)? mem[1324] : 
                         (N119)? mem[1388] : 
                         (N121)? mem[1452] : 
                         (N123)? mem[1516] : 
                         (N125)? mem[1580] : 
                         (N127)? mem[1644] : 
                         (N129)? mem[1708] : 
                         (N131)? mem[1772] : 
                         (N133)? mem[1836] : 
                         (N135)? mem[1900] : 
                         (N137)? mem[1964] : 
                         (N139)? mem[2028] : 1'b0;
  assign r1_data_o[43] = (N108)? mem[43] : 
                         (N110)? mem[107] : 
                         (N112)? mem[171] : 
                         (N114)? mem[235] : 
                         (N116)? mem[299] : 
                         (N118)? mem[363] : 
                         (N120)? mem[427] : 
                         (N122)? mem[491] : 
                         (N124)? mem[555] : 
                         (N126)? mem[619] : 
                         (N128)? mem[683] : 
                         (N130)? mem[747] : 
                         (N132)? mem[811] : 
                         (N134)? mem[875] : 
                         (N136)? mem[939] : 
                         (N138)? mem[1003] : 
                         (N109)? mem[1067] : 
                         (N111)? mem[1131] : 
                         (N113)? mem[1195] : 
                         (N115)? mem[1259] : 
                         (N117)? mem[1323] : 
                         (N119)? mem[1387] : 
                         (N121)? mem[1451] : 
                         (N123)? mem[1515] : 
                         (N125)? mem[1579] : 
                         (N127)? mem[1643] : 
                         (N129)? mem[1707] : 
                         (N131)? mem[1771] : 
                         (N133)? mem[1835] : 
                         (N135)? mem[1899] : 
                         (N137)? mem[1963] : 
                         (N139)? mem[2027] : 1'b0;
  assign r1_data_o[42] = (N108)? mem[42] : 
                         (N110)? mem[106] : 
                         (N112)? mem[170] : 
                         (N114)? mem[234] : 
                         (N116)? mem[298] : 
                         (N118)? mem[362] : 
                         (N120)? mem[426] : 
                         (N122)? mem[490] : 
                         (N124)? mem[554] : 
                         (N126)? mem[618] : 
                         (N128)? mem[682] : 
                         (N130)? mem[746] : 
                         (N132)? mem[810] : 
                         (N134)? mem[874] : 
                         (N136)? mem[938] : 
                         (N138)? mem[1002] : 
                         (N109)? mem[1066] : 
                         (N111)? mem[1130] : 
                         (N113)? mem[1194] : 
                         (N115)? mem[1258] : 
                         (N117)? mem[1322] : 
                         (N119)? mem[1386] : 
                         (N121)? mem[1450] : 
                         (N123)? mem[1514] : 
                         (N125)? mem[1578] : 
                         (N127)? mem[1642] : 
                         (N129)? mem[1706] : 
                         (N131)? mem[1770] : 
                         (N133)? mem[1834] : 
                         (N135)? mem[1898] : 
                         (N137)? mem[1962] : 
                         (N139)? mem[2026] : 1'b0;
  assign r1_data_o[41] = (N108)? mem[41] : 
                         (N110)? mem[105] : 
                         (N112)? mem[169] : 
                         (N114)? mem[233] : 
                         (N116)? mem[297] : 
                         (N118)? mem[361] : 
                         (N120)? mem[425] : 
                         (N122)? mem[489] : 
                         (N124)? mem[553] : 
                         (N126)? mem[617] : 
                         (N128)? mem[681] : 
                         (N130)? mem[745] : 
                         (N132)? mem[809] : 
                         (N134)? mem[873] : 
                         (N136)? mem[937] : 
                         (N138)? mem[1001] : 
                         (N109)? mem[1065] : 
                         (N111)? mem[1129] : 
                         (N113)? mem[1193] : 
                         (N115)? mem[1257] : 
                         (N117)? mem[1321] : 
                         (N119)? mem[1385] : 
                         (N121)? mem[1449] : 
                         (N123)? mem[1513] : 
                         (N125)? mem[1577] : 
                         (N127)? mem[1641] : 
                         (N129)? mem[1705] : 
                         (N131)? mem[1769] : 
                         (N133)? mem[1833] : 
                         (N135)? mem[1897] : 
                         (N137)? mem[1961] : 
                         (N139)? mem[2025] : 1'b0;
  assign r1_data_o[40] = (N108)? mem[40] : 
                         (N110)? mem[104] : 
                         (N112)? mem[168] : 
                         (N114)? mem[232] : 
                         (N116)? mem[296] : 
                         (N118)? mem[360] : 
                         (N120)? mem[424] : 
                         (N122)? mem[488] : 
                         (N124)? mem[552] : 
                         (N126)? mem[616] : 
                         (N128)? mem[680] : 
                         (N130)? mem[744] : 
                         (N132)? mem[808] : 
                         (N134)? mem[872] : 
                         (N136)? mem[936] : 
                         (N138)? mem[1000] : 
                         (N109)? mem[1064] : 
                         (N111)? mem[1128] : 
                         (N113)? mem[1192] : 
                         (N115)? mem[1256] : 
                         (N117)? mem[1320] : 
                         (N119)? mem[1384] : 
                         (N121)? mem[1448] : 
                         (N123)? mem[1512] : 
                         (N125)? mem[1576] : 
                         (N127)? mem[1640] : 
                         (N129)? mem[1704] : 
                         (N131)? mem[1768] : 
                         (N133)? mem[1832] : 
                         (N135)? mem[1896] : 
                         (N137)? mem[1960] : 
                         (N139)? mem[2024] : 1'b0;
  assign r1_data_o[39] = (N108)? mem[39] : 
                         (N110)? mem[103] : 
                         (N112)? mem[167] : 
                         (N114)? mem[231] : 
                         (N116)? mem[295] : 
                         (N118)? mem[359] : 
                         (N120)? mem[423] : 
                         (N122)? mem[487] : 
                         (N124)? mem[551] : 
                         (N126)? mem[615] : 
                         (N128)? mem[679] : 
                         (N130)? mem[743] : 
                         (N132)? mem[807] : 
                         (N134)? mem[871] : 
                         (N136)? mem[935] : 
                         (N138)? mem[999] : 
                         (N109)? mem[1063] : 
                         (N111)? mem[1127] : 
                         (N113)? mem[1191] : 
                         (N115)? mem[1255] : 
                         (N117)? mem[1319] : 
                         (N119)? mem[1383] : 
                         (N121)? mem[1447] : 
                         (N123)? mem[1511] : 
                         (N125)? mem[1575] : 
                         (N127)? mem[1639] : 
                         (N129)? mem[1703] : 
                         (N131)? mem[1767] : 
                         (N133)? mem[1831] : 
                         (N135)? mem[1895] : 
                         (N137)? mem[1959] : 
                         (N139)? mem[2023] : 1'b0;
  assign r1_data_o[38] = (N108)? mem[38] : 
                         (N110)? mem[102] : 
                         (N112)? mem[166] : 
                         (N114)? mem[230] : 
                         (N116)? mem[294] : 
                         (N118)? mem[358] : 
                         (N120)? mem[422] : 
                         (N122)? mem[486] : 
                         (N124)? mem[550] : 
                         (N126)? mem[614] : 
                         (N128)? mem[678] : 
                         (N130)? mem[742] : 
                         (N132)? mem[806] : 
                         (N134)? mem[870] : 
                         (N136)? mem[934] : 
                         (N138)? mem[998] : 
                         (N109)? mem[1062] : 
                         (N111)? mem[1126] : 
                         (N113)? mem[1190] : 
                         (N115)? mem[1254] : 
                         (N117)? mem[1318] : 
                         (N119)? mem[1382] : 
                         (N121)? mem[1446] : 
                         (N123)? mem[1510] : 
                         (N125)? mem[1574] : 
                         (N127)? mem[1638] : 
                         (N129)? mem[1702] : 
                         (N131)? mem[1766] : 
                         (N133)? mem[1830] : 
                         (N135)? mem[1894] : 
                         (N137)? mem[1958] : 
                         (N139)? mem[2022] : 1'b0;
  assign r1_data_o[37] = (N108)? mem[37] : 
                         (N110)? mem[101] : 
                         (N112)? mem[165] : 
                         (N114)? mem[229] : 
                         (N116)? mem[293] : 
                         (N118)? mem[357] : 
                         (N120)? mem[421] : 
                         (N122)? mem[485] : 
                         (N124)? mem[549] : 
                         (N126)? mem[613] : 
                         (N128)? mem[677] : 
                         (N130)? mem[741] : 
                         (N132)? mem[805] : 
                         (N134)? mem[869] : 
                         (N136)? mem[933] : 
                         (N138)? mem[997] : 
                         (N109)? mem[1061] : 
                         (N111)? mem[1125] : 
                         (N113)? mem[1189] : 
                         (N115)? mem[1253] : 
                         (N117)? mem[1317] : 
                         (N119)? mem[1381] : 
                         (N121)? mem[1445] : 
                         (N123)? mem[1509] : 
                         (N125)? mem[1573] : 
                         (N127)? mem[1637] : 
                         (N129)? mem[1701] : 
                         (N131)? mem[1765] : 
                         (N133)? mem[1829] : 
                         (N135)? mem[1893] : 
                         (N137)? mem[1957] : 
                         (N139)? mem[2021] : 1'b0;
  assign r1_data_o[36] = (N108)? mem[36] : 
                         (N110)? mem[100] : 
                         (N112)? mem[164] : 
                         (N114)? mem[228] : 
                         (N116)? mem[292] : 
                         (N118)? mem[356] : 
                         (N120)? mem[420] : 
                         (N122)? mem[484] : 
                         (N124)? mem[548] : 
                         (N126)? mem[612] : 
                         (N128)? mem[676] : 
                         (N130)? mem[740] : 
                         (N132)? mem[804] : 
                         (N134)? mem[868] : 
                         (N136)? mem[932] : 
                         (N138)? mem[996] : 
                         (N109)? mem[1060] : 
                         (N111)? mem[1124] : 
                         (N113)? mem[1188] : 
                         (N115)? mem[1252] : 
                         (N117)? mem[1316] : 
                         (N119)? mem[1380] : 
                         (N121)? mem[1444] : 
                         (N123)? mem[1508] : 
                         (N125)? mem[1572] : 
                         (N127)? mem[1636] : 
                         (N129)? mem[1700] : 
                         (N131)? mem[1764] : 
                         (N133)? mem[1828] : 
                         (N135)? mem[1892] : 
                         (N137)? mem[1956] : 
                         (N139)? mem[2020] : 1'b0;
  assign r1_data_o[35] = (N108)? mem[35] : 
                         (N110)? mem[99] : 
                         (N112)? mem[163] : 
                         (N114)? mem[227] : 
                         (N116)? mem[291] : 
                         (N118)? mem[355] : 
                         (N120)? mem[419] : 
                         (N122)? mem[483] : 
                         (N124)? mem[547] : 
                         (N126)? mem[611] : 
                         (N128)? mem[675] : 
                         (N130)? mem[739] : 
                         (N132)? mem[803] : 
                         (N134)? mem[867] : 
                         (N136)? mem[931] : 
                         (N138)? mem[995] : 
                         (N109)? mem[1059] : 
                         (N111)? mem[1123] : 
                         (N113)? mem[1187] : 
                         (N115)? mem[1251] : 
                         (N117)? mem[1315] : 
                         (N119)? mem[1379] : 
                         (N121)? mem[1443] : 
                         (N123)? mem[1507] : 
                         (N125)? mem[1571] : 
                         (N127)? mem[1635] : 
                         (N129)? mem[1699] : 
                         (N131)? mem[1763] : 
                         (N133)? mem[1827] : 
                         (N135)? mem[1891] : 
                         (N137)? mem[1955] : 
                         (N139)? mem[2019] : 1'b0;
  assign r1_data_o[34] = (N108)? mem[34] : 
                         (N110)? mem[98] : 
                         (N112)? mem[162] : 
                         (N114)? mem[226] : 
                         (N116)? mem[290] : 
                         (N118)? mem[354] : 
                         (N120)? mem[418] : 
                         (N122)? mem[482] : 
                         (N124)? mem[546] : 
                         (N126)? mem[610] : 
                         (N128)? mem[674] : 
                         (N130)? mem[738] : 
                         (N132)? mem[802] : 
                         (N134)? mem[866] : 
                         (N136)? mem[930] : 
                         (N138)? mem[994] : 
                         (N109)? mem[1058] : 
                         (N111)? mem[1122] : 
                         (N113)? mem[1186] : 
                         (N115)? mem[1250] : 
                         (N117)? mem[1314] : 
                         (N119)? mem[1378] : 
                         (N121)? mem[1442] : 
                         (N123)? mem[1506] : 
                         (N125)? mem[1570] : 
                         (N127)? mem[1634] : 
                         (N129)? mem[1698] : 
                         (N131)? mem[1762] : 
                         (N133)? mem[1826] : 
                         (N135)? mem[1890] : 
                         (N137)? mem[1954] : 
                         (N139)? mem[2018] : 1'b0;
  assign r1_data_o[33] = (N108)? mem[33] : 
                         (N110)? mem[97] : 
                         (N112)? mem[161] : 
                         (N114)? mem[225] : 
                         (N116)? mem[289] : 
                         (N118)? mem[353] : 
                         (N120)? mem[417] : 
                         (N122)? mem[481] : 
                         (N124)? mem[545] : 
                         (N126)? mem[609] : 
                         (N128)? mem[673] : 
                         (N130)? mem[737] : 
                         (N132)? mem[801] : 
                         (N134)? mem[865] : 
                         (N136)? mem[929] : 
                         (N138)? mem[993] : 
                         (N109)? mem[1057] : 
                         (N111)? mem[1121] : 
                         (N113)? mem[1185] : 
                         (N115)? mem[1249] : 
                         (N117)? mem[1313] : 
                         (N119)? mem[1377] : 
                         (N121)? mem[1441] : 
                         (N123)? mem[1505] : 
                         (N125)? mem[1569] : 
                         (N127)? mem[1633] : 
                         (N129)? mem[1697] : 
                         (N131)? mem[1761] : 
                         (N133)? mem[1825] : 
                         (N135)? mem[1889] : 
                         (N137)? mem[1953] : 
                         (N139)? mem[2017] : 1'b0;
  assign r1_data_o[32] = (N108)? mem[32] : 
                         (N110)? mem[96] : 
                         (N112)? mem[160] : 
                         (N114)? mem[224] : 
                         (N116)? mem[288] : 
                         (N118)? mem[352] : 
                         (N120)? mem[416] : 
                         (N122)? mem[480] : 
                         (N124)? mem[544] : 
                         (N126)? mem[608] : 
                         (N128)? mem[672] : 
                         (N130)? mem[736] : 
                         (N132)? mem[800] : 
                         (N134)? mem[864] : 
                         (N136)? mem[928] : 
                         (N138)? mem[992] : 
                         (N109)? mem[1056] : 
                         (N111)? mem[1120] : 
                         (N113)? mem[1184] : 
                         (N115)? mem[1248] : 
                         (N117)? mem[1312] : 
                         (N119)? mem[1376] : 
                         (N121)? mem[1440] : 
                         (N123)? mem[1504] : 
                         (N125)? mem[1568] : 
                         (N127)? mem[1632] : 
                         (N129)? mem[1696] : 
                         (N131)? mem[1760] : 
                         (N133)? mem[1824] : 
                         (N135)? mem[1888] : 
                         (N137)? mem[1952] : 
                         (N139)? mem[2016] : 1'b0;
  assign r1_data_o[31] = (N108)? mem[31] : 
                         (N110)? mem[95] : 
                         (N112)? mem[159] : 
                         (N114)? mem[223] : 
                         (N116)? mem[287] : 
                         (N118)? mem[351] : 
                         (N120)? mem[415] : 
                         (N122)? mem[479] : 
                         (N124)? mem[543] : 
                         (N126)? mem[607] : 
                         (N128)? mem[671] : 
                         (N130)? mem[735] : 
                         (N132)? mem[799] : 
                         (N134)? mem[863] : 
                         (N136)? mem[927] : 
                         (N138)? mem[991] : 
                         (N109)? mem[1055] : 
                         (N111)? mem[1119] : 
                         (N113)? mem[1183] : 
                         (N115)? mem[1247] : 
                         (N117)? mem[1311] : 
                         (N119)? mem[1375] : 
                         (N121)? mem[1439] : 
                         (N123)? mem[1503] : 
                         (N125)? mem[1567] : 
                         (N127)? mem[1631] : 
                         (N129)? mem[1695] : 
                         (N131)? mem[1759] : 
                         (N133)? mem[1823] : 
                         (N135)? mem[1887] : 
                         (N137)? mem[1951] : 
                         (N139)? mem[2015] : 1'b0;
  assign r1_data_o[30] = (N108)? mem[30] : 
                         (N110)? mem[94] : 
                         (N112)? mem[158] : 
                         (N114)? mem[222] : 
                         (N116)? mem[286] : 
                         (N118)? mem[350] : 
                         (N120)? mem[414] : 
                         (N122)? mem[478] : 
                         (N124)? mem[542] : 
                         (N126)? mem[606] : 
                         (N128)? mem[670] : 
                         (N130)? mem[734] : 
                         (N132)? mem[798] : 
                         (N134)? mem[862] : 
                         (N136)? mem[926] : 
                         (N138)? mem[990] : 
                         (N109)? mem[1054] : 
                         (N111)? mem[1118] : 
                         (N113)? mem[1182] : 
                         (N115)? mem[1246] : 
                         (N117)? mem[1310] : 
                         (N119)? mem[1374] : 
                         (N121)? mem[1438] : 
                         (N123)? mem[1502] : 
                         (N125)? mem[1566] : 
                         (N127)? mem[1630] : 
                         (N129)? mem[1694] : 
                         (N131)? mem[1758] : 
                         (N133)? mem[1822] : 
                         (N135)? mem[1886] : 
                         (N137)? mem[1950] : 
                         (N139)? mem[2014] : 1'b0;
  assign r1_data_o[29] = (N108)? mem[29] : 
                         (N110)? mem[93] : 
                         (N112)? mem[157] : 
                         (N114)? mem[221] : 
                         (N116)? mem[285] : 
                         (N118)? mem[349] : 
                         (N120)? mem[413] : 
                         (N122)? mem[477] : 
                         (N124)? mem[541] : 
                         (N126)? mem[605] : 
                         (N128)? mem[669] : 
                         (N130)? mem[733] : 
                         (N132)? mem[797] : 
                         (N134)? mem[861] : 
                         (N136)? mem[925] : 
                         (N138)? mem[989] : 
                         (N109)? mem[1053] : 
                         (N111)? mem[1117] : 
                         (N113)? mem[1181] : 
                         (N115)? mem[1245] : 
                         (N117)? mem[1309] : 
                         (N119)? mem[1373] : 
                         (N121)? mem[1437] : 
                         (N123)? mem[1501] : 
                         (N125)? mem[1565] : 
                         (N127)? mem[1629] : 
                         (N129)? mem[1693] : 
                         (N131)? mem[1757] : 
                         (N133)? mem[1821] : 
                         (N135)? mem[1885] : 
                         (N137)? mem[1949] : 
                         (N139)? mem[2013] : 1'b0;
  assign r1_data_o[28] = (N108)? mem[28] : 
                         (N110)? mem[92] : 
                         (N112)? mem[156] : 
                         (N114)? mem[220] : 
                         (N116)? mem[284] : 
                         (N118)? mem[348] : 
                         (N120)? mem[412] : 
                         (N122)? mem[476] : 
                         (N124)? mem[540] : 
                         (N126)? mem[604] : 
                         (N128)? mem[668] : 
                         (N130)? mem[732] : 
                         (N132)? mem[796] : 
                         (N134)? mem[860] : 
                         (N136)? mem[924] : 
                         (N138)? mem[988] : 
                         (N109)? mem[1052] : 
                         (N111)? mem[1116] : 
                         (N113)? mem[1180] : 
                         (N115)? mem[1244] : 
                         (N117)? mem[1308] : 
                         (N119)? mem[1372] : 
                         (N121)? mem[1436] : 
                         (N123)? mem[1500] : 
                         (N125)? mem[1564] : 
                         (N127)? mem[1628] : 
                         (N129)? mem[1692] : 
                         (N131)? mem[1756] : 
                         (N133)? mem[1820] : 
                         (N135)? mem[1884] : 
                         (N137)? mem[1948] : 
                         (N139)? mem[2012] : 1'b0;
  assign r1_data_o[27] = (N108)? mem[27] : 
                         (N110)? mem[91] : 
                         (N112)? mem[155] : 
                         (N114)? mem[219] : 
                         (N116)? mem[283] : 
                         (N118)? mem[347] : 
                         (N120)? mem[411] : 
                         (N122)? mem[475] : 
                         (N124)? mem[539] : 
                         (N126)? mem[603] : 
                         (N128)? mem[667] : 
                         (N130)? mem[731] : 
                         (N132)? mem[795] : 
                         (N134)? mem[859] : 
                         (N136)? mem[923] : 
                         (N138)? mem[987] : 
                         (N109)? mem[1051] : 
                         (N111)? mem[1115] : 
                         (N113)? mem[1179] : 
                         (N115)? mem[1243] : 
                         (N117)? mem[1307] : 
                         (N119)? mem[1371] : 
                         (N121)? mem[1435] : 
                         (N123)? mem[1499] : 
                         (N125)? mem[1563] : 
                         (N127)? mem[1627] : 
                         (N129)? mem[1691] : 
                         (N131)? mem[1755] : 
                         (N133)? mem[1819] : 
                         (N135)? mem[1883] : 
                         (N137)? mem[1947] : 
                         (N139)? mem[2011] : 1'b0;
  assign r1_data_o[26] = (N108)? mem[26] : 
                         (N110)? mem[90] : 
                         (N112)? mem[154] : 
                         (N114)? mem[218] : 
                         (N116)? mem[282] : 
                         (N118)? mem[346] : 
                         (N120)? mem[410] : 
                         (N122)? mem[474] : 
                         (N124)? mem[538] : 
                         (N126)? mem[602] : 
                         (N128)? mem[666] : 
                         (N130)? mem[730] : 
                         (N132)? mem[794] : 
                         (N134)? mem[858] : 
                         (N136)? mem[922] : 
                         (N138)? mem[986] : 
                         (N109)? mem[1050] : 
                         (N111)? mem[1114] : 
                         (N113)? mem[1178] : 
                         (N115)? mem[1242] : 
                         (N117)? mem[1306] : 
                         (N119)? mem[1370] : 
                         (N121)? mem[1434] : 
                         (N123)? mem[1498] : 
                         (N125)? mem[1562] : 
                         (N127)? mem[1626] : 
                         (N129)? mem[1690] : 
                         (N131)? mem[1754] : 
                         (N133)? mem[1818] : 
                         (N135)? mem[1882] : 
                         (N137)? mem[1946] : 
                         (N139)? mem[2010] : 1'b0;
  assign r1_data_o[25] = (N108)? mem[25] : 
                         (N110)? mem[89] : 
                         (N112)? mem[153] : 
                         (N114)? mem[217] : 
                         (N116)? mem[281] : 
                         (N118)? mem[345] : 
                         (N120)? mem[409] : 
                         (N122)? mem[473] : 
                         (N124)? mem[537] : 
                         (N126)? mem[601] : 
                         (N128)? mem[665] : 
                         (N130)? mem[729] : 
                         (N132)? mem[793] : 
                         (N134)? mem[857] : 
                         (N136)? mem[921] : 
                         (N138)? mem[985] : 
                         (N109)? mem[1049] : 
                         (N111)? mem[1113] : 
                         (N113)? mem[1177] : 
                         (N115)? mem[1241] : 
                         (N117)? mem[1305] : 
                         (N119)? mem[1369] : 
                         (N121)? mem[1433] : 
                         (N123)? mem[1497] : 
                         (N125)? mem[1561] : 
                         (N127)? mem[1625] : 
                         (N129)? mem[1689] : 
                         (N131)? mem[1753] : 
                         (N133)? mem[1817] : 
                         (N135)? mem[1881] : 
                         (N137)? mem[1945] : 
                         (N139)? mem[2009] : 1'b0;
  assign r1_data_o[24] = (N108)? mem[24] : 
                         (N110)? mem[88] : 
                         (N112)? mem[152] : 
                         (N114)? mem[216] : 
                         (N116)? mem[280] : 
                         (N118)? mem[344] : 
                         (N120)? mem[408] : 
                         (N122)? mem[472] : 
                         (N124)? mem[536] : 
                         (N126)? mem[600] : 
                         (N128)? mem[664] : 
                         (N130)? mem[728] : 
                         (N132)? mem[792] : 
                         (N134)? mem[856] : 
                         (N136)? mem[920] : 
                         (N138)? mem[984] : 
                         (N109)? mem[1048] : 
                         (N111)? mem[1112] : 
                         (N113)? mem[1176] : 
                         (N115)? mem[1240] : 
                         (N117)? mem[1304] : 
                         (N119)? mem[1368] : 
                         (N121)? mem[1432] : 
                         (N123)? mem[1496] : 
                         (N125)? mem[1560] : 
                         (N127)? mem[1624] : 
                         (N129)? mem[1688] : 
                         (N131)? mem[1752] : 
                         (N133)? mem[1816] : 
                         (N135)? mem[1880] : 
                         (N137)? mem[1944] : 
                         (N139)? mem[2008] : 1'b0;
  assign r1_data_o[23] = (N108)? mem[23] : 
                         (N110)? mem[87] : 
                         (N112)? mem[151] : 
                         (N114)? mem[215] : 
                         (N116)? mem[279] : 
                         (N118)? mem[343] : 
                         (N120)? mem[407] : 
                         (N122)? mem[471] : 
                         (N124)? mem[535] : 
                         (N126)? mem[599] : 
                         (N128)? mem[663] : 
                         (N130)? mem[727] : 
                         (N132)? mem[791] : 
                         (N134)? mem[855] : 
                         (N136)? mem[919] : 
                         (N138)? mem[983] : 
                         (N109)? mem[1047] : 
                         (N111)? mem[1111] : 
                         (N113)? mem[1175] : 
                         (N115)? mem[1239] : 
                         (N117)? mem[1303] : 
                         (N119)? mem[1367] : 
                         (N121)? mem[1431] : 
                         (N123)? mem[1495] : 
                         (N125)? mem[1559] : 
                         (N127)? mem[1623] : 
                         (N129)? mem[1687] : 
                         (N131)? mem[1751] : 
                         (N133)? mem[1815] : 
                         (N135)? mem[1879] : 
                         (N137)? mem[1943] : 
                         (N139)? mem[2007] : 1'b0;
  assign r1_data_o[22] = (N108)? mem[22] : 
                         (N110)? mem[86] : 
                         (N112)? mem[150] : 
                         (N114)? mem[214] : 
                         (N116)? mem[278] : 
                         (N118)? mem[342] : 
                         (N120)? mem[406] : 
                         (N122)? mem[470] : 
                         (N124)? mem[534] : 
                         (N126)? mem[598] : 
                         (N128)? mem[662] : 
                         (N130)? mem[726] : 
                         (N132)? mem[790] : 
                         (N134)? mem[854] : 
                         (N136)? mem[918] : 
                         (N138)? mem[982] : 
                         (N109)? mem[1046] : 
                         (N111)? mem[1110] : 
                         (N113)? mem[1174] : 
                         (N115)? mem[1238] : 
                         (N117)? mem[1302] : 
                         (N119)? mem[1366] : 
                         (N121)? mem[1430] : 
                         (N123)? mem[1494] : 
                         (N125)? mem[1558] : 
                         (N127)? mem[1622] : 
                         (N129)? mem[1686] : 
                         (N131)? mem[1750] : 
                         (N133)? mem[1814] : 
                         (N135)? mem[1878] : 
                         (N137)? mem[1942] : 
                         (N139)? mem[2006] : 1'b0;
  assign r1_data_o[21] = (N108)? mem[21] : 
                         (N110)? mem[85] : 
                         (N112)? mem[149] : 
                         (N114)? mem[213] : 
                         (N116)? mem[277] : 
                         (N118)? mem[341] : 
                         (N120)? mem[405] : 
                         (N122)? mem[469] : 
                         (N124)? mem[533] : 
                         (N126)? mem[597] : 
                         (N128)? mem[661] : 
                         (N130)? mem[725] : 
                         (N132)? mem[789] : 
                         (N134)? mem[853] : 
                         (N136)? mem[917] : 
                         (N138)? mem[981] : 
                         (N109)? mem[1045] : 
                         (N111)? mem[1109] : 
                         (N113)? mem[1173] : 
                         (N115)? mem[1237] : 
                         (N117)? mem[1301] : 
                         (N119)? mem[1365] : 
                         (N121)? mem[1429] : 
                         (N123)? mem[1493] : 
                         (N125)? mem[1557] : 
                         (N127)? mem[1621] : 
                         (N129)? mem[1685] : 
                         (N131)? mem[1749] : 
                         (N133)? mem[1813] : 
                         (N135)? mem[1877] : 
                         (N137)? mem[1941] : 
                         (N139)? mem[2005] : 1'b0;
  assign r1_data_o[20] = (N108)? mem[20] : 
                         (N110)? mem[84] : 
                         (N112)? mem[148] : 
                         (N114)? mem[212] : 
                         (N116)? mem[276] : 
                         (N118)? mem[340] : 
                         (N120)? mem[404] : 
                         (N122)? mem[468] : 
                         (N124)? mem[532] : 
                         (N126)? mem[596] : 
                         (N128)? mem[660] : 
                         (N130)? mem[724] : 
                         (N132)? mem[788] : 
                         (N134)? mem[852] : 
                         (N136)? mem[916] : 
                         (N138)? mem[980] : 
                         (N109)? mem[1044] : 
                         (N111)? mem[1108] : 
                         (N113)? mem[1172] : 
                         (N115)? mem[1236] : 
                         (N117)? mem[1300] : 
                         (N119)? mem[1364] : 
                         (N121)? mem[1428] : 
                         (N123)? mem[1492] : 
                         (N125)? mem[1556] : 
                         (N127)? mem[1620] : 
                         (N129)? mem[1684] : 
                         (N131)? mem[1748] : 
                         (N133)? mem[1812] : 
                         (N135)? mem[1876] : 
                         (N137)? mem[1940] : 
                         (N139)? mem[2004] : 1'b0;
  assign r1_data_o[19] = (N108)? mem[19] : 
                         (N110)? mem[83] : 
                         (N112)? mem[147] : 
                         (N114)? mem[211] : 
                         (N116)? mem[275] : 
                         (N118)? mem[339] : 
                         (N120)? mem[403] : 
                         (N122)? mem[467] : 
                         (N124)? mem[531] : 
                         (N126)? mem[595] : 
                         (N128)? mem[659] : 
                         (N130)? mem[723] : 
                         (N132)? mem[787] : 
                         (N134)? mem[851] : 
                         (N136)? mem[915] : 
                         (N138)? mem[979] : 
                         (N109)? mem[1043] : 
                         (N111)? mem[1107] : 
                         (N113)? mem[1171] : 
                         (N115)? mem[1235] : 
                         (N117)? mem[1299] : 
                         (N119)? mem[1363] : 
                         (N121)? mem[1427] : 
                         (N123)? mem[1491] : 
                         (N125)? mem[1555] : 
                         (N127)? mem[1619] : 
                         (N129)? mem[1683] : 
                         (N131)? mem[1747] : 
                         (N133)? mem[1811] : 
                         (N135)? mem[1875] : 
                         (N137)? mem[1939] : 
                         (N139)? mem[2003] : 1'b0;
  assign r1_data_o[18] = (N108)? mem[18] : 
                         (N110)? mem[82] : 
                         (N112)? mem[146] : 
                         (N114)? mem[210] : 
                         (N116)? mem[274] : 
                         (N118)? mem[338] : 
                         (N120)? mem[402] : 
                         (N122)? mem[466] : 
                         (N124)? mem[530] : 
                         (N126)? mem[594] : 
                         (N128)? mem[658] : 
                         (N130)? mem[722] : 
                         (N132)? mem[786] : 
                         (N134)? mem[850] : 
                         (N136)? mem[914] : 
                         (N138)? mem[978] : 
                         (N109)? mem[1042] : 
                         (N111)? mem[1106] : 
                         (N113)? mem[1170] : 
                         (N115)? mem[1234] : 
                         (N117)? mem[1298] : 
                         (N119)? mem[1362] : 
                         (N121)? mem[1426] : 
                         (N123)? mem[1490] : 
                         (N125)? mem[1554] : 
                         (N127)? mem[1618] : 
                         (N129)? mem[1682] : 
                         (N131)? mem[1746] : 
                         (N133)? mem[1810] : 
                         (N135)? mem[1874] : 
                         (N137)? mem[1938] : 
                         (N139)? mem[2002] : 1'b0;
  assign r1_data_o[17] = (N108)? mem[17] : 
                         (N110)? mem[81] : 
                         (N112)? mem[145] : 
                         (N114)? mem[209] : 
                         (N116)? mem[273] : 
                         (N118)? mem[337] : 
                         (N120)? mem[401] : 
                         (N122)? mem[465] : 
                         (N124)? mem[529] : 
                         (N126)? mem[593] : 
                         (N128)? mem[657] : 
                         (N130)? mem[721] : 
                         (N132)? mem[785] : 
                         (N134)? mem[849] : 
                         (N136)? mem[913] : 
                         (N138)? mem[977] : 
                         (N109)? mem[1041] : 
                         (N111)? mem[1105] : 
                         (N113)? mem[1169] : 
                         (N115)? mem[1233] : 
                         (N117)? mem[1297] : 
                         (N119)? mem[1361] : 
                         (N121)? mem[1425] : 
                         (N123)? mem[1489] : 
                         (N125)? mem[1553] : 
                         (N127)? mem[1617] : 
                         (N129)? mem[1681] : 
                         (N131)? mem[1745] : 
                         (N133)? mem[1809] : 
                         (N135)? mem[1873] : 
                         (N137)? mem[1937] : 
                         (N139)? mem[2001] : 1'b0;
  assign r1_data_o[16] = (N108)? mem[16] : 
                         (N110)? mem[80] : 
                         (N112)? mem[144] : 
                         (N114)? mem[208] : 
                         (N116)? mem[272] : 
                         (N118)? mem[336] : 
                         (N120)? mem[400] : 
                         (N122)? mem[464] : 
                         (N124)? mem[528] : 
                         (N126)? mem[592] : 
                         (N128)? mem[656] : 
                         (N130)? mem[720] : 
                         (N132)? mem[784] : 
                         (N134)? mem[848] : 
                         (N136)? mem[912] : 
                         (N138)? mem[976] : 
                         (N109)? mem[1040] : 
                         (N111)? mem[1104] : 
                         (N113)? mem[1168] : 
                         (N115)? mem[1232] : 
                         (N117)? mem[1296] : 
                         (N119)? mem[1360] : 
                         (N121)? mem[1424] : 
                         (N123)? mem[1488] : 
                         (N125)? mem[1552] : 
                         (N127)? mem[1616] : 
                         (N129)? mem[1680] : 
                         (N131)? mem[1744] : 
                         (N133)? mem[1808] : 
                         (N135)? mem[1872] : 
                         (N137)? mem[1936] : 
                         (N139)? mem[2000] : 1'b0;
  assign r1_data_o[15] = (N108)? mem[15] : 
                         (N110)? mem[79] : 
                         (N112)? mem[143] : 
                         (N114)? mem[207] : 
                         (N116)? mem[271] : 
                         (N118)? mem[335] : 
                         (N120)? mem[399] : 
                         (N122)? mem[463] : 
                         (N124)? mem[527] : 
                         (N126)? mem[591] : 
                         (N128)? mem[655] : 
                         (N130)? mem[719] : 
                         (N132)? mem[783] : 
                         (N134)? mem[847] : 
                         (N136)? mem[911] : 
                         (N138)? mem[975] : 
                         (N109)? mem[1039] : 
                         (N111)? mem[1103] : 
                         (N113)? mem[1167] : 
                         (N115)? mem[1231] : 
                         (N117)? mem[1295] : 
                         (N119)? mem[1359] : 
                         (N121)? mem[1423] : 
                         (N123)? mem[1487] : 
                         (N125)? mem[1551] : 
                         (N127)? mem[1615] : 
                         (N129)? mem[1679] : 
                         (N131)? mem[1743] : 
                         (N133)? mem[1807] : 
                         (N135)? mem[1871] : 
                         (N137)? mem[1935] : 
                         (N139)? mem[1999] : 1'b0;
  assign r1_data_o[14] = (N108)? mem[14] : 
                         (N110)? mem[78] : 
                         (N112)? mem[142] : 
                         (N114)? mem[206] : 
                         (N116)? mem[270] : 
                         (N118)? mem[334] : 
                         (N120)? mem[398] : 
                         (N122)? mem[462] : 
                         (N124)? mem[526] : 
                         (N126)? mem[590] : 
                         (N128)? mem[654] : 
                         (N130)? mem[718] : 
                         (N132)? mem[782] : 
                         (N134)? mem[846] : 
                         (N136)? mem[910] : 
                         (N138)? mem[974] : 
                         (N109)? mem[1038] : 
                         (N111)? mem[1102] : 
                         (N113)? mem[1166] : 
                         (N115)? mem[1230] : 
                         (N117)? mem[1294] : 
                         (N119)? mem[1358] : 
                         (N121)? mem[1422] : 
                         (N123)? mem[1486] : 
                         (N125)? mem[1550] : 
                         (N127)? mem[1614] : 
                         (N129)? mem[1678] : 
                         (N131)? mem[1742] : 
                         (N133)? mem[1806] : 
                         (N135)? mem[1870] : 
                         (N137)? mem[1934] : 
                         (N139)? mem[1998] : 1'b0;
  assign r1_data_o[13] = (N108)? mem[13] : 
                         (N110)? mem[77] : 
                         (N112)? mem[141] : 
                         (N114)? mem[205] : 
                         (N116)? mem[269] : 
                         (N118)? mem[333] : 
                         (N120)? mem[397] : 
                         (N122)? mem[461] : 
                         (N124)? mem[525] : 
                         (N126)? mem[589] : 
                         (N128)? mem[653] : 
                         (N130)? mem[717] : 
                         (N132)? mem[781] : 
                         (N134)? mem[845] : 
                         (N136)? mem[909] : 
                         (N138)? mem[973] : 
                         (N109)? mem[1037] : 
                         (N111)? mem[1101] : 
                         (N113)? mem[1165] : 
                         (N115)? mem[1229] : 
                         (N117)? mem[1293] : 
                         (N119)? mem[1357] : 
                         (N121)? mem[1421] : 
                         (N123)? mem[1485] : 
                         (N125)? mem[1549] : 
                         (N127)? mem[1613] : 
                         (N129)? mem[1677] : 
                         (N131)? mem[1741] : 
                         (N133)? mem[1805] : 
                         (N135)? mem[1869] : 
                         (N137)? mem[1933] : 
                         (N139)? mem[1997] : 1'b0;
  assign r1_data_o[12] = (N108)? mem[12] : 
                         (N110)? mem[76] : 
                         (N112)? mem[140] : 
                         (N114)? mem[204] : 
                         (N116)? mem[268] : 
                         (N118)? mem[332] : 
                         (N120)? mem[396] : 
                         (N122)? mem[460] : 
                         (N124)? mem[524] : 
                         (N126)? mem[588] : 
                         (N128)? mem[652] : 
                         (N130)? mem[716] : 
                         (N132)? mem[780] : 
                         (N134)? mem[844] : 
                         (N136)? mem[908] : 
                         (N138)? mem[972] : 
                         (N109)? mem[1036] : 
                         (N111)? mem[1100] : 
                         (N113)? mem[1164] : 
                         (N115)? mem[1228] : 
                         (N117)? mem[1292] : 
                         (N119)? mem[1356] : 
                         (N121)? mem[1420] : 
                         (N123)? mem[1484] : 
                         (N125)? mem[1548] : 
                         (N127)? mem[1612] : 
                         (N129)? mem[1676] : 
                         (N131)? mem[1740] : 
                         (N133)? mem[1804] : 
                         (N135)? mem[1868] : 
                         (N137)? mem[1932] : 
                         (N139)? mem[1996] : 1'b0;
  assign r1_data_o[11] = (N108)? mem[11] : 
                         (N110)? mem[75] : 
                         (N112)? mem[139] : 
                         (N114)? mem[203] : 
                         (N116)? mem[267] : 
                         (N118)? mem[331] : 
                         (N120)? mem[395] : 
                         (N122)? mem[459] : 
                         (N124)? mem[523] : 
                         (N126)? mem[587] : 
                         (N128)? mem[651] : 
                         (N130)? mem[715] : 
                         (N132)? mem[779] : 
                         (N134)? mem[843] : 
                         (N136)? mem[907] : 
                         (N138)? mem[971] : 
                         (N109)? mem[1035] : 
                         (N111)? mem[1099] : 
                         (N113)? mem[1163] : 
                         (N115)? mem[1227] : 
                         (N117)? mem[1291] : 
                         (N119)? mem[1355] : 
                         (N121)? mem[1419] : 
                         (N123)? mem[1483] : 
                         (N125)? mem[1547] : 
                         (N127)? mem[1611] : 
                         (N129)? mem[1675] : 
                         (N131)? mem[1739] : 
                         (N133)? mem[1803] : 
                         (N135)? mem[1867] : 
                         (N137)? mem[1931] : 
                         (N139)? mem[1995] : 1'b0;
  assign r1_data_o[10] = (N108)? mem[10] : 
                         (N110)? mem[74] : 
                         (N112)? mem[138] : 
                         (N114)? mem[202] : 
                         (N116)? mem[266] : 
                         (N118)? mem[330] : 
                         (N120)? mem[394] : 
                         (N122)? mem[458] : 
                         (N124)? mem[522] : 
                         (N126)? mem[586] : 
                         (N128)? mem[650] : 
                         (N130)? mem[714] : 
                         (N132)? mem[778] : 
                         (N134)? mem[842] : 
                         (N136)? mem[906] : 
                         (N138)? mem[970] : 
                         (N109)? mem[1034] : 
                         (N111)? mem[1098] : 
                         (N113)? mem[1162] : 
                         (N115)? mem[1226] : 
                         (N117)? mem[1290] : 
                         (N119)? mem[1354] : 
                         (N121)? mem[1418] : 
                         (N123)? mem[1482] : 
                         (N125)? mem[1546] : 
                         (N127)? mem[1610] : 
                         (N129)? mem[1674] : 
                         (N131)? mem[1738] : 
                         (N133)? mem[1802] : 
                         (N135)? mem[1866] : 
                         (N137)? mem[1930] : 
                         (N139)? mem[1994] : 1'b0;
  assign r1_data_o[9] = (N108)? mem[9] : 
                        (N110)? mem[73] : 
                        (N112)? mem[137] : 
                        (N114)? mem[201] : 
                        (N116)? mem[265] : 
                        (N118)? mem[329] : 
                        (N120)? mem[393] : 
                        (N122)? mem[457] : 
                        (N124)? mem[521] : 
                        (N126)? mem[585] : 
                        (N128)? mem[649] : 
                        (N130)? mem[713] : 
                        (N132)? mem[777] : 
                        (N134)? mem[841] : 
                        (N136)? mem[905] : 
                        (N138)? mem[969] : 
                        (N109)? mem[1033] : 
                        (N111)? mem[1097] : 
                        (N113)? mem[1161] : 
                        (N115)? mem[1225] : 
                        (N117)? mem[1289] : 
                        (N119)? mem[1353] : 
                        (N121)? mem[1417] : 
                        (N123)? mem[1481] : 
                        (N125)? mem[1545] : 
                        (N127)? mem[1609] : 
                        (N129)? mem[1673] : 
                        (N131)? mem[1737] : 
                        (N133)? mem[1801] : 
                        (N135)? mem[1865] : 
                        (N137)? mem[1929] : 
                        (N139)? mem[1993] : 1'b0;
  assign r1_data_o[8] = (N108)? mem[8] : 
                        (N110)? mem[72] : 
                        (N112)? mem[136] : 
                        (N114)? mem[200] : 
                        (N116)? mem[264] : 
                        (N118)? mem[328] : 
                        (N120)? mem[392] : 
                        (N122)? mem[456] : 
                        (N124)? mem[520] : 
                        (N126)? mem[584] : 
                        (N128)? mem[648] : 
                        (N130)? mem[712] : 
                        (N132)? mem[776] : 
                        (N134)? mem[840] : 
                        (N136)? mem[904] : 
                        (N138)? mem[968] : 
                        (N109)? mem[1032] : 
                        (N111)? mem[1096] : 
                        (N113)? mem[1160] : 
                        (N115)? mem[1224] : 
                        (N117)? mem[1288] : 
                        (N119)? mem[1352] : 
                        (N121)? mem[1416] : 
                        (N123)? mem[1480] : 
                        (N125)? mem[1544] : 
                        (N127)? mem[1608] : 
                        (N129)? mem[1672] : 
                        (N131)? mem[1736] : 
                        (N133)? mem[1800] : 
                        (N135)? mem[1864] : 
                        (N137)? mem[1928] : 
                        (N139)? mem[1992] : 1'b0;
  assign r1_data_o[7] = (N108)? mem[7] : 
                        (N110)? mem[71] : 
                        (N112)? mem[135] : 
                        (N114)? mem[199] : 
                        (N116)? mem[263] : 
                        (N118)? mem[327] : 
                        (N120)? mem[391] : 
                        (N122)? mem[455] : 
                        (N124)? mem[519] : 
                        (N126)? mem[583] : 
                        (N128)? mem[647] : 
                        (N130)? mem[711] : 
                        (N132)? mem[775] : 
                        (N134)? mem[839] : 
                        (N136)? mem[903] : 
                        (N138)? mem[967] : 
                        (N109)? mem[1031] : 
                        (N111)? mem[1095] : 
                        (N113)? mem[1159] : 
                        (N115)? mem[1223] : 
                        (N117)? mem[1287] : 
                        (N119)? mem[1351] : 
                        (N121)? mem[1415] : 
                        (N123)? mem[1479] : 
                        (N125)? mem[1543] : 
                        (N127)? mem[1607] : 
                        (N129)? mem[1671] : 
                        (N131)? mem[1735] : 
                        (N133)? mem[1799] : 
                        (N135)? mem[1863] : 
                        (N137)? mem[1927] : 
                        (N139)? mem[1991] : 1'b0;
  assign r1_data_o[6] = (N108)? mem[6] : 
                        (N110)? mem[70] : 
                        (N112)? mem[134] : 
                        (N114)? mem[198] : 
                        (N116)? mem[262] : 
                        (N118)? mem[326] : 
                        (N120)? mem[390] : 
                        (N122)? mem[454] : 
                        (N124)? mem[518] : 
                        (N126)? mem[582] : 
                        (N128)? mem[646] : 
                        (N130)? mem[710] : 
                        (N132)? mem[774] : 
                        (N134)? mem[838] : 
                        (N136)? mem[902] : 
                        (N138)? mem[966] : 
                        (N109)? mem[1030] : 
                        (N111)? mem[1094] : 
                        (N113)? mem[1158] : 
                        (N115)? mem[1222] : 
                        (N117)? mem[1286] : 
                        (N119)? mem[1350] : 
                        (N121)? mem[1414] : 
                        (N123)? mem[1478] : 
                        (N125)? mem[1542] : 
                        (N127)? mem[1606] : 
                        (N129)? mem[1670] : 
                        (N131)? mem[1734] : 
                        (N133)? mem[1798] : 
                        (N135)? mem[1862] : 
                        (N137)? mem[1926] : 
                        (N139)? mem[1990] : 1'b0;
  assign r1_data_o[5] = (N108)? mem[5] : 
                        (N110)? mem[69] : 
                        (N112)? mem[133] : 
                        (N114)? mem[197] : 
                        (N116)? mem[261] : 
                        (N118)? mem[325] : 
                        (N120)? mem[389] : 
                        (N122)? mem[453] : 
                        (N124)? mem[517] : 
                        (N126)? mem[581] : 
                        (N128)? mem[645] : 
                        (N130)? mem[709] : 
                        (N132)? mem[773] : 
                        (N134)? mem[837] : 
                        (N136)? mem[901] : 
                        (N138)? mem[965] : 
                        (N109)? mem[1029] : 
                        (N111)? mem[1093] : 
                        (N113)? mem[1157] : 
                        (N115)? mem[1221] : 
                        (N117)? mem[1285] : 
                        (N119)? mem[1349] : 
                        (N121)? mem[1413] : 
                        (N123)? mem[1477] : 
                        (N125)? mem[1541] : 
                        (N127)? mem[1605] : 
                        (N129)? mem[1669] : 
                        (N131)? mem[1733] : 
                        (N133)? mem[1797] : 
                        (N135)? mem[1861] : 
                        (N137)? mem[1925] : 
                        (N139)? mem[1989] : 1'b0;
  assign r1_data_o[4] = (N108)? mem[4] : 
                        (N110)? mem[68] : 
                        (N112)? mem[132] : 
                        (N114)? mem[196] : 
                        (N116)? mem[260] : 
                        (N118)? mem[324] : 
                        (N120)? mem[388] : 
                        (N122)? mem[452] : 
                        (N124)? mem[516] : 
                        (N126)? mem[580] : 
                        (N128)? mem[644] : 
                        (N130)? mem[708] : 
                        (N132)? mem[772] : 
                        (N134)? mem[836] : 
                        (N136)? mem[900] : 
                        (N138)? mem[964] : 
                        (N109)? mem[1028] : 
                        (N111)? mem[1092] : 
                        (N113)? mem[1156] : 
                        (N115)? mem[1220] : 
                        (N117)? mem[1284] : 
                        (N119)? mem[1348] : 
                        (N121)? mem[1412] : 
                        (N123)? mem[1476] : 
                        (N125)? mem[1540] : 
                        (N127)? mem[1604] : 
                        (N129)? mem[1668] : 
                        (N131)? mem[1732] : 
                        (N133)? mem[1796] : 
                        (N135)? mem[1860] : 
                        (N137)? mem[1924] : 
                        (N139)? mem[1988] : 1'b0;
  assign r1_data_o[3] = (N108)? mem[3] : 
                        (N110)? mem[67] : 
                        (N112)? mem[131] : 
                        (N114)? mem[195] : 
                        (N116)? mem[259] : 
                        (N118)? mem[323] : 
                        (N120)? mem[387] : 
                        (N122)? mem[451] : 
                        (N124)? mem[515] : 
                        (N126)? mem[579] : 
                        (N128)? mem[643] : 
                        (N130)? mem[707] : 
                        (N132)? mem[771] : 
                        (N134)? mem[835] : 
                        (N136)? mem[899] : 
                        (N138)? mem[963] : 
                        (N109)? mem[1027] : 
                        (N111)? mem[1091] : 
                        (N113)? mem[1155] : 
                        (N115)? mem[1219] : 
                        (N117)? mem[1283] : 
                        (N119)? mem[1347] : 
                        (N121)? mem[1411] : 
                        (N123)? mem[1475] : 
                        (N125)? mem[1539] : 
                        (N127)? mem[1603] : 
                        (N129)? mem[1667] : 
                        (N131)? mem[1731] : 
                        (N133)? mem[1795] : 
                        (N135)? mem[1859] : 
                        (N137)? mem[1923] : 
                        (N139)? mem[1987] : 1'b0;
  assign r1_data_o[2] = (N108)? mem[2] : 
                        (N110)? mem[66] : 
                        (N112)? mem[130] : 
                        (N114)? mem[194] : 
                        (N116)? mem[258] : 
                        (N118)? mem[322] : 
                        (N120)? mem[386] : 
                        (N122)? mem[450] : 
                        (N124)? mem[514] : 
                        (N126)? mem[578] : 
                        (N128)? mem[642] : 
                        (N130)? mem[706] : 
                        (N132)? mem[770] : 
                        (N134)? mem[834] : 
                        (N136)? mem[898] : 
                        (N138)? mem[962] : 
                        (N109)? mem[1026] : 
                        (N111)? mem[1090] : 
                        (N113)? mem[1154] : 
                        (N115)? mem[1218] : 
                        (N117)? mem[1282] : 
                        (N119)? mem[1346] : 
                        (N121)? mem[1410] : 
                        (N123)? mem[1474] : 
                        (N125)? mem[1538] : 
                        (N127)? mem[1602] : 
                        (N129)? mem[1666] : 
                        (N131)? mem[1730] : 
                        (N133)? mem[1794] : 
                        (N135)? mem[1858] : 
                        (N137)? mem[1922] : 
                        (N139)? mem[1986] : 1'b0;
  assign r1_data_o[1] = (N108)? mem[1] : 
                        (N110)? mem[65] : 
                        (N112)? mem[129] : 
                        (N114)? mem[193] : 
                        (N116)? mem[257] : 
                        (N118)? mem[321] : 
                        (N120)? mem[385] : 
                        (N122)? mem[449] : 
                        (N124)? mem[513] : 
                        (N126)? mem[577] : 
                        (N128)? mem[641] : 
                        (N130)? mem[705] : 
                        (N132)? mem[769] : 
                        (N134)? mem[833] : 
                        (N136)? mem[897] : 
                        (N138)? mem[961] : 
                        (N109)? mem[1025] : 
                        (N111)? mem[1089] : 
                        (N113)? mem[1153] : 
                        (N115)? mem[1217] : 
                        (N117)? mem[1281] : 
                        (N119)? mem[1345] : 
                        (N121)? mem[1409] : 
                        (N123)? mem[1473] : 
                        (N125)? mem[1537] : 
                        (N127)? mem[1601] : 
                        (N129)? mem[1665] : 
                        (N131)? mem[1729] : 
                        (N133)? mem[1793] : 
                        (N135)? mem[1857] : 
                        (N137)? mem[1921] : 
                        (N139)? mem[1985] : 1'b0;
  assign r1_data_o[0] = (N108)? mem[0] : 
                        (N110)? mem[64] : 
                        (N112)? mem[128] : 
                        (N114)? mem[192] : 
                        (N116)? mem[256] : 
                        (N118)? mem[320] : 
                        (N120)? mem[384] : 
                        (N122)? mem[448] : 
                        (N124)? mem[512] : 
                        (N126)? mem[576] : 
                        (N128)? mem[640] : 
                        (N130)? mem[704] : 
                        (N132)? mem[768] : 
                        (N134)? mem[832] : 
                        (N136)? mem[896] : 
                        (N138)? mem[960] : 
                        (N109)? mem[1024] : 
                        (N111)? mem[1088] : 
                        (N113)? mem[1152] : 
                        (N115)? mem[1216] : 
                        (N117)? mem[1280] : 
                        (N119)? mem[1344] : 
                        (N121)? mem[1408] : 
                        (N123)? mem[1472] : 
                        (N125)? mem[1536] : 
                        (N127)? mem[1600] : 
                        (N129)? mem[1664] : 
                        (N131)? mem[1728] : 
                        (N133)? mem[1792] : 
                        (N135)? mem[1856] : 
                        (N137)? mem[1920] : 
                        (N139)? mem[1984] : 1'b0;
  assign N205 = w_addr_i[3] & w_addr_i[4];
  assign N206 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N207 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N208 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N209 = ~w_addr_i[2];
  assign N210 = w_addr_i[0] & w_addr_i[1];
  assign N211 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N212 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N213 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N214 = w_addr_i[2] & N210;
  assign N215 = w_addr_i[2] & N211;
  assign N216 = w_addr_i[2] & N212;
  assign N217 = w_addr_i[2] & N213;
  assign N218 = N209 & N210;
  assign N219 = N209 & N211;
  assign N220 = N209 & N212;
  assign N221 = N209 & N213;
  assign N172 = N205 & N214;
  assign N171 = N205 & N215;
  assign N170 = N205 & N216;
  assign N169 = N205 & N217;
  assign N168 = N205 & N218;
  assign N167 = N205 & N219;
  assign N166 = N205 & N220;
  assign N165 = N205 & N221;
  assign N164 = N206 & N214;
  assign N163 = N206 & N215;
  assign N162 = N206 & N216;
  assign N161 = N206 & N217;
  assign N160 = N206 & N218;
  assign N159 = N206 & N219;
  assign N158 = N206 & N220;
  assign N157 = N206 & N221;
  assign N156 = N207 & N214;
  assign N155 = N207 & N215;
  assign N154 = N207 & N216;
  assign N153 = N207 & N217;
  assign N152 = N207 & N218;
  assign N151 = N207 & N219;
  assign N150 = N207 & N220;
  assign N149 = N207 & N221;
  assign N148 = N208 & N214;
  assign N147 = N208 & N215;
  assign N146 = N208 & N216;
  assign N145 = N208 & N217;
  assign N144 = N208 & N218;
  assign N143 = N208 & N219;
  assign N142 = N208 & N220;
  assign N141 = N208 & N221;
  assign { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173 } = (N8)? { N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141 } : 
                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N140;
  assign N10 = ~r0_addr_r[0];
  assign N11 = ~r0_addr_r[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r0_addr_r[1];
  assign N14 = r0_addr_r[0] & N11;
  assign N15 = r0_addr_r[0] & r0_addr_r[1];
  assign N16 = ~r0_addr_r[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r0_addr_r[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r0_addr_r[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r0_addr_r[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r0_addr_r[2];
  assign N25 = ~r0_addr_r[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r0_addr_r[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r0_addr_r[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r0_addr_r[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r0_addr_r[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r0_addr_r[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r0_addr_r[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r0_addr_r[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r0_addr_r[3];
  assign N42 = ~r0_addr_r[4];
  assign N43 = N26 & N42;
  assign N44 = N26 & r0_addr_r[4];
  assign N45 = N28 & N42;
  assign N46 = N28 & r0_addr_r[4];
  assign N47 = N30 & N42;
  assign N48 = N30 & r0_addr_r[4];
  assign N49 = N32 & N42;
  assign N50 = N32 & r0_addr_r[4];
  assign N51 = N34 & N42;
  assign N52 = N34 & r0_addr_r[4];
  assign N53 = N36 & N42;
  assign N54 = N36 & r0_addr_r[4];
  assign N55 = N38 & N42;
  assign N56 = N38 & r0_addr_r[4];
  assign N57 = N40 & N42;
  assign N58 = N40 & r0_addr_r[4];
  assign N59 = N27 & N42;
  assign N60 = N27 & r0_addr_r[4];
  assign N61 = N29 & N42;
  assign N62 = N29 & r0_addr_r[4];
  assign N63 = N31 & N42;
  assign N64 = N31 & r0_addr_r[4];
  assign N65 = N33 & N42;
  assign N66 = N33 & r0_addr_r[4];
  assign N67 = N35 & N42;
  assign N68 = N35 & r0_addr_r[4];
  assign N69 = N37 & N42;
  assign N70 = N37 & r0_addr_r[4];
  assign N71 = N39 & N42;
  assign N72 = N39 & r0_addr_r[4];
  assign N73 = N41 & N42;
  assign N74 = N41 & r0_addr_r[4];
  assign N75 = ~r1_addr_r[0];
  assign N76 = ~r1_addr_r[1];
  assign N77 = N75 & N76;
  assign N78 = N75 & r1_addr_r[1];
  assign N79 = r1_addr_r[0] & N76;
  assign N80 = r1_addr_r[0] & r1_addr_r[1];
  assign N81 = ~r1_addr_r[2];
  assign N82 = N77 & N81;
  assign N83 = N77 & r1_addr_r[2];
  assign N84 = N79 & N81;
  assign N85 = N79 & r1_addr_r[2];
  assign N86 = N78 & N81;
  assign N87 = N78 & r1_addr_r[2];
  assign N88 = N80 & N81;
  assign N89 = N80 & r1_addr_r[2];
  assign N90 = ~r1_addr_r[3];
  assign N91 = N82 & N90;
  assign N92 = N82 & r1_addr_r[3];
  assign N93 = N84 & N90;
  assign N94 = N84 & r1_addr_r[3];
  assign N95 = N86 & N90;
  assign N96 = N86 & r1_addr_r[3];
  assign N97 = N88 & N90;
  assign N98 = N88 & r1_addr_r[3];
  assign N99 = N83 & N90;
  assign N100 = N83 & r1_addr_r[3];
  assign N101 = N85 & N90;
  assign N102 = N85 & r1_addr_r[3];
  assign N103 = N87 & N90;
  assign N104 = N87 & r1_addr_r[3];
  assign N105 = N89 & N90;
  assign N106 = N89 & r1_addr_r[3];
  assign N107 = ~r1_addr_r[4];
  assign N108 = N91 & N107;
  assign N109 = N91 & r1_addr_r[4];
  assign N110 = N93 & N107;
  assign N111 = N93 & r1_addr_r[4];
  assign N112 = N95 & N107;
  assign N113 = N95 & r1_addr_r[4];
  assign N114 = N97 & N107;
  assign N115 = N97 & r1_addr_r[4];
  assign N116 = N99 & N107;
  assign N117 = N99 & r1_addr_r[4];
  assign N118 = N101 & N107;
  assign N119 = N101 & r1_addr_r[4];
  assign N120 = N103 & N107;
  assign N121 = N103 & r1_addr_r[4];
  assign N122 = N105 & N107;
  assign N123 = N105 & r1_addr_r[4];
  assign N124 = N92 & N107;
  assign N125 = N92 & r1_addr_r[4];
  assign N126 = N94 & N107;
  assign N127 = N94 & r1_addr_r[4];
  assign N128 = N96 & N107;
  assign N129 = N96 & r1_addr_r[4];
  assign N130 = N98 & N107;
  assign N131 = N98 & r1_addr_r[4];
  assign N132 = N100 & N107;
  assign N133 = N100 & r1_addr_r[4];
  assign N134 = N102 & N107;
  assign N135 = N102 & r1_addr_r[4];
  assign N136 = N104 & N107;
  assign N137 = N104 & r1_addr_r[4];
  assign N138 = N106 & N107;
  assign N139 = N106 & r1_addr_r[4];
  assign N140 = ~w_v_i;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { r0_addr_r[4:0] } <= { r0_addr_i[4:0] };
      { r1_addr_r[4:0] } <= { r1_addr_i[4:0] };
    end 
    if(N204) begin
      { mem[2047:1984] } <= { w_data_i[63:0] };
    end 
    if(N203) begin
      { mem[1983:1920] } <= { w_data_i[63:0] };
    end 
    if(N202) begin
      { mem[1919:1856] } <= { w_data_i[63:0] };
    end 
    if(N201) begin
      { mem[1855:1792] } <= { w_data_i[63:0] };
    end 
    if(N200) begin
      { mem[1791:1728] } <= { w_data_i[63:0] };
    end 
    if(N199) begin
      { mem[1727:1664] } <= { w_data_i[63:0] };
    end 
    if(N198) begin
      { mem[1663:1600] } <= { w_data_i[63:0] };
    end 
    if(N197) begin
      { mem[1599:1536] } <= { w_data_i[63:0] };
    end 
    if(N196) begin
      { mem[1535:1472] } <= { w_data_i[63:0] };
    end 
    if(N195) begin
      { mem[1471:1408] } <= { w_data_i[63:0] };
    end 
    if(N194) begin
      { mem[1407:1344] } <= { w_data_i[63:0] };
    end 
    if(N193) begin
      { mem[1343:1280] } <= { w_data_i[63:0] };
    end 
    if(N192) begin
      { mem[1279:1216] } <= { w_data_i[63:0] };
    end 
    if(N191) begin
      { mem[1215:1152] } <= { w_data_i[63:0] };
    end 
    if(N190) begin
      { mem[1151:1088] } <= { w_data_i[63:0] };
    end 
    if(N189) begin
      { mem[1087:1024] } <= { w_data_i[63:0] };
    end 
    if(N188) begin
      { mem[1023:960] } <= { w_data_i[63:0] };
    end 
    if(N187) begin
      { mem[959:896] } <= { w_data_i[63:0] };
    end 
    if(N186) begin
      { mem[895:832] } <= { w_data_i[63:0] };
    end 
    if(N185) begin
      { mem[831:768] } <= { w_data_i[63:0] };
    end 
    if(N184) begin
      { mem[767:704] } <= { w_data_i[63:0] };
    end 
    if(N183) begin
      { mem[703:640] } <= { w_data_i[63:0] };
    end 
    if(N182) begin
      { mem[639:576] } <= { w_data_i[63:0] };
    end 
    if(N181) begin
      { mem[575:512] } <= { w_data_i[63:0] };
    end 
    if(N180) begin
      { mem[511:448] } <= { w_data_i[63:0] };
    end 
    if(N179) begin
      { mem[447:384] } <= { w_data_i[63:0] };
    end 
    if(N178) begin
      { mem[383:320] } <= { w_data_i[63:0] };
    end 
    if(N177) begin
      { mem[319:256] } <= { w_data_i[63:0] };
    end 
    if(N176) begin
      { mem[255:192] } <= { w_data_i[63:0] };
    end 
    if(N175) begin
      { mem[191:128] } <= { w_data_i[63:0] };
    end 
    if(N174) begin
      { mem[127:64] } <= { w_data_i[63:0] };
    end 
    if(N173) begin
      { mem[63:0] } <= { w_data_i[63:0] };
    end 
  end


endmodule



module bsg_mem_2r1w_sync_width_p64_els_p32_read_write_same_addr_p1
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r0_v_i,
  r0_addr_i,
  r0_data_o,
  r1_v_i,
  r1_addr_i,
  r1_data_o
);

  input [4:0] w_addr_i;
  input [63:0] w_data_i;
  input [4:0] r0_addr_i;
  output [63:0] r0_data_o;
  input [4:0] r1_addr_i;
  output [63:0] r1_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r0_v_i;
  input r1_v_i;
  wire [63:0] r0_data_o,r1_data_o;

  bsg_mem_2r1w_sync_synth_width_p64_els_p32_read_write_same_addr_p1_harden_p0
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r0_v_i(r0_v_i),
    .r0_addr_i(r0_addr_i),
    .r0_data_o(r0_data_o),
    .r1_v_i(r1_v_i),
    .r1_addr_i(r1_addr_i),
    .r1_data_o(r1_data_o)
  );


endmodule



module bsg_dff_en_width_p5
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [4:0] data_i;
  output [4:0] data_o;
  input clk_i;
  input en_i;
  reg [4:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[4:0] } <= { data_i[4:0] };
    end 
  end


endmodule



module bp_be_regfile
(
  clk_i,
  reset_i,
  issue_v_i,
  dispatch_v_i,
  rd_w_v_i,
  rd_addr_i,
  rd_data_i,
  rs1_r_v_i,
  rs1_addr_i,
  rs1_data_o,
  rs2_r_v_i,
  rs2_addr_i,
  rs2_data_o
);

  input [4:0] rd_addr_i;
  input [63:0] rd_data_i;
  input [4:0] rs1_addr_i;
  output [63:0] rs1_data_o;
  input [4:0] rs2_addr_i;
  output [63:0] rs2_data_o;
  input clk_i;
  input reset_i;
  input issue_v_i;
  input dispatch_v_i;
  input rd_w_v_i;
  input rs1_r_v_i;
  input rs2_r_v_i;
  wire [63:0] rs1_data_o,rs2_data_o,rs1_reg_data,rs2_reg_data;
  wire N0,N1,N2,N3,N4,N5,N6,N7,rs1_read_v,rs2_read_v,rs1_issue_v,rs2_issue_v,N8,N9,N10,
  N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;
  wire [4:0] rs1_reread_addr,rs2_reread_addr,rs1_addr_r,rs2_addr_r;

  bsg_mem_2r1w_sync_width_p64_els_p32_read_write_same_addr_p1
  rf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(rd_w_v_i),
    .w_addr_i(rd_addr_i),
    .w_data_i(rd_data_i),
    .r0_v_i(rs1_read_v),
    .r0_addr_i(rs1_reread_addr),
    .r0_data_o(rs1_reg_data),
    .r1_v_i(rs2_read_v),
    .r1_addr_i(rs2_reread_addr),
    .r1_data_o(rs2_reg_data)
  );


  bsg_dff_en_width_p5
  rs1_addr
  (
    .clk_i(clk_i),
    .data_i(rs1_addr_i),
    .en_i(rs1_issue_v),
    .data_o(rs1_addr_r)
  );


  bsg_dff_en_width_p5
  rs2_addr
  (
    .clk_i(clk_i),
    .data_i(rs2_addr_i),
    .en_i(rs2_issue_v),
    .data_o(rs2_addr_r)
  );

  assign N12 = rs1_addr_r[3] | rs1_addr_r[4];
  assign N13 = rs1_addr_r[2] | N12;
  assign N14 = rs1_addr_r[1] | N13;
  assign N15 = rs1_addr_r[0] | N14;
  assign N16 = ~N15;
  assign N17 = rs2_addr_r[3] | rs2_addr_r[4];
  assign N18 = rs2_addr_r[2] | N17;
  assign N19 = rs2_addr_r[1] | N18;
  assign N20 = rs2_addr_r[0] | N19;
  assign N21 = ~N20;
  assign rs1_reread_addr = (N0)? rs1_addr_i : 
                           (N1)? rs1_addr_r : 1'b0;
  assign N0 = N9;
  assign N1 = N8;
  assign rs2_reread_addr = (N2)? rs2_addr_i : 
                           (N3)? rs2_addr_r : 1'b0;
  assign N2 = N11;
  assign N3 = N10;
  assign rs1_data_o = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N5)? rs1_reg_data : 1'b0;
  assign N4 = N16;
  assign N5 = N15;
  assign rs2_data_o = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N7)? rs2_reg_data : 1'b0;
  assign N6 = N21;
  assign N7 = N20;
  assign rs1_issue_v = issue_v_i & rs1_r_v_i;
  assign rs2_issue_v = issue_v_i & rs2_r_v_i;
  assign rs1_read_v = rs1_issue_v | N22;
  assign N22 = ~dispatch_v_i;
  assign rs2_read_v = rs2_issue_v | N22;
  assign N8 = ~rs1_issue_v;
  assign N9 = rs1_issue_v;
  assign N10 = ~rs2_issue_v;
  assign N11 = rs2_issue_v;

endmodule



module bsg_dff_reset_en_width_p221
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [220:0] data_i;
  output [220:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228;
  reg [220:0] data_o;
  assign { N7, N5, N3 } = (N0)? { 1'b1, 1'b1, 1'b1 } : 
                          (N228)? { 1'b1, 1'b1, 1'b1 } : 
                          (N2)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = reset_i;
  assign { N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N6, N4 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N228)? data_i : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N227 = ~reset_i;
  assign N228 = en_i & N227;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[220:122], data_o[0:0] } <= { N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N4 };
    end 
    if(N5) begin
      { data_o[121:23], data_o[1:1] } <= { N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N6 };
    end 
    if(N7) begin
      { data_o[22:2] } <= { N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8 };
    end 
  end


endmodule



module bp_be_instr_decoder
(
  instr_i,
  fe_nop_v_i,
  be_nop_v_i,
  me_nop_v_i,
  decode_o,
  illegal_instr_o
);

  input [31:0] instr_i;
  output [42:0] decode_o;
  input fe_nop_v_i;
  input be_nop_v_i;
  input me_nop_v_i;
  output illegal_instr_o;
  wire [42:0] decode_o;
  wire illegal_instr_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,
  N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,
  N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,
  N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,
  N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,
  N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,
  N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,
  N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,
  N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
  N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,
  N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,
  N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,
  N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,
  N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,
  N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
  N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,
  N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,
  N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,
  N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
  N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,
  N370,N371,N372;
  assign decode_o[26] = 1'b0;
  assign decode_o[27] = 1'b0;
  assign decode_o[28] = 1'b0;
  assign decode_o[32] = 1'b0;
  assign decode_o[34] = 1'b0;
  assign decode_o[36] = 1'b0;
  assign N54 = instr_i[1] & instr_i[0];
  assign N56 = instr_i[6] | N339;
  assign N57 = N340 | instr_i[3];
  assign N58 = N56 | N57;
  assign N59 = N58 | instr_i[2];
  assign N60 = N340 | N341;
  assign N61 = N56 | N60;
  assign N62 = N61 | instr_i[2];
  assign N64 = instr_i[6] | instr_i[5];
  assign N65 = N64 | N57;
  assign N66 = N65 | instr_i[2];
  assign N67 = N64 | N60;
  assign N68 = N67 | instr_i[2];
  assign N70 = N58 | N86;
  assign N72 = N65 | N86;
  assign N74 = N85 | N339;
  assign N75 = instr_i[4] | N341;
  assign N76 = N74 | N75;
  assign N77 = N76 | N86;
  assign N79 = instr_i[4] | instr_i[3];
  assign N80 = N74 | N79;
  assign N81 = N80 | N86;
  assign N83 = N80 | instr_i[2];
  assign N87 = N85 & N339;
  assign N88 = N340 & N341;
  assign N89 = N87 & N88;
  assign N90 = N89 & N86;
  assign N91 = N56 | N79;
  assign N92 = N91 | instr_i[2];
  assign N94 = N64 | N75;
  assign N95 = N94 | N86;
  assign N97 = N74 | N57;
  assign N98 = N97 | instr_i[2];
  assign N100 = instr_i[6] & instr_i[4];
  assign N101 = N100 & instr_i[2];
  assign N102 = N100 & instr_i[3];
  assign N103 = instr_i[4] & instr_i[3];
  assign N104 = N103 & instr_i[2];
  assign N105 = N85 & instr_i[5];
  assign N106 = N340 & instr_i[2];
  assign N107 = N105 & N106;
  assign N108 = N85 & N340;
  assign N109 = N341 & instr_i[2];
  assign N110 = N108 & N109;
  assign N111 = N339 & N340;
  assign N112 = N111 & N109;
  assign N113 = N340 & instr_i[3];
  assign N114 = N113 & N86;
  assign N115 = instr_i[6] & N339;
  assign N123 = N117 & N118;
  assign N124 = N119 & N120;
  assign N125 = N121 & N122;
  assign N126 = instr_i[4] & N86;
  assign N127 = N123 & N124;
  assign N128 = N125 & N105;
  assign N129 = N126 & N54;
  assign N130 = N127 & N128;
  assign N131 = N130 & N129;
  assign N133 = N154 & N285;
  assign N134 = N133 & N341;
  assign N135 = N133 & instr_i[3];
  assign N137 = N166 & N285;
  assign N138 = N137 & N341;
  assign N139 = N137 & instr_i[3];
  assign N141 = N154 & N286;
  assign N142 = N141 & N341;
  assign N143 = N141 & instr_i[3];
  assign N145 = N159 & N286;
  assign N146 = N145 & N341;
  assign N147 = N145 & instr_i[3];
  assign N149 = N172 & N286;
  assign N150 = N149 & N341;
  assign N151 = N149 & instr_i[3];
  assign N154 = N153 & N251;
  assign N155 = N154 & N287;
  assign N156 = N155 & N341;
  assign N157 = N154 & N288;
  assign N158 = N157 & N341;
  assign N159 = N153 & instr_i[14];
  assign N160 = N159 & N285;
  assign N161 = N160 & N341;
  assign N162 = N159 & N287;
  assign N163 = N162 & N341;
  assign N164 = N159 & N288;
  assign N165 = N164 & N341;
  assign N166 = instr_i[30] & N251;
  assign N167 = N166 & instr_i[12];
  assign N168 = instr_i[14] & N284;
  assign N169 = N168 & instr_i[3];
  assign N170 = instr_i[13] & instr_i[3];
  assign N171 = instr_i[30] & instr_i[13];
  assign N172 = instr_i[30] & instr_i[14];
  assign N173 = N172 & N284;
  assign N185 = N87 & N126;
  assign N186 = N185 & N54;
  assign N188 = N242 & N216;
  assign N189 = N284 & instr_i[3];
  assign N190 = N242 & N189;
  assign N192 = N205 & N242;
  assign N193 = N198 & N192;
  assign N194 = N193 & N218;
  assign N195 = N193 & N210;
  assign N197 = N117 & N153;
  assign N198 = N197 & N204;
  assign N199 = N198 & N207;
  assign N200 = N199 & N218;
  assign N201 = N199 & N210;
  assign N203 = N117 & instr_i[30];
  assign N204 = N118 & N119;
  assign N205 = N120 & N121;
  assign N206 = N203 & N204;
  assign N207 = N205 & N245;
  assign N208 = N206 & N207;
  assign N209 = N208 & N218;
  assign N210 = instr_i[12] & instr_i[3];
  assign N211 = N208 & N210;
  assign N213 = N252 & N216;
  assign N214 = N252 & N218;
  assign N215 = N245 & N216;
  assign N216 = N284 & N341;
  assign N217 = N248 & N216;
  assign N218 = instr_i[12] & N341;
  assign N219 = N248 & N218;
  assign N238 = instr_i[2] | N342;
  assign N239 = N238 | N343;
  assign N240 = N80 | N239;
  assign N242 = N251 & N283;
  assign N243 = N242 & N284;
  assign N244 = N242 & instr_i[12];
  assign N245 = instr_i[14] & N283;
  assign N246 = N245 & N284;
  assign N247 = N245 & instr_i[12];
  assign N248 = instr_i[14] & instr_i[13];
  assign N249 = N248 & N284;
  assign N250 = N248 & instr_i[12];
  assign N252 = N251 & instr_i[13];
  assign N263 = N64 | N79;
  assign N264 = N263 | N239;
  assign N266 = N252 & N284;
  assign N267 = N252 & instr_i[12];
  assign N276 = N251 & N85;
  assign N277 = instr_i[5] & N340;
  assign N278 = N341 & N86;
  assign N279 = N276 & N277;
  assign N280 = N278 & N54;
  assign N281 = N279 & N280;
  assign N285 = N283 & N284;
  assign N286 = N283 & instr_i[12];
  assign N287 = instr_i[13] & N284;
  assign N288 = instr_i[13] & instr_i[12];
  assign N296 = N117 | N153;
  assign N297 = N118 | N119;
  assign N298 = instr_i[27] | instr_i[26];
  assign N299 = instr_i[25] | N294;
  assign N300 = instr_i[23] | N295;
  assign N301 = instr_i[21] | instr_i[20];
  assign N302 = N296 | N297;
  assign N303 = N298 | N299;
  assign N304 = N300 | N301;
  assign N305 = N302 | N303;
  assign N306 = N305 | N304;
  assign N339 = ~instr_i[5];
  assign N340 = ~instr_i[4];
  assign N341 = ~instr_i[3];
  assign N342 = ~instr_i[1];
  assign N343 = ~instr_i[0];
  assign N344 = N339 | instr_i[6];
  assign N345 = N340 | N344;
  assign N346 = N341 | N345;
  assign N347 = instr_i[2] | N346;
  assign N348 = N342 | N347;
  assign N349 = N343 | N348;
  assign N350 = ~N349;
  assign N351 = instr_i[5] | instr_i[6];
  assign N352 = N340 | N351;
  assign N353 = N341 | N352;
  assign N354 = instr_i[2] | N353;
  assign N355 = N342 | N354;
  assign N356 = N343 | N355;
  assign N357 = ~N356;
  assign { N178, N177, N176, N175 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N1)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N2)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                      (N3)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                      (N4)? { 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                      (N5)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N6)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                      (N7)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                      (N8)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                      (N9)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                      (N10)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N136;
  assign N1 = N140;
  assign N2 = N144;
  assign N3 = N148;
  assign N4 = N152;
  assign N5 = N156;
  assign N6 = N158;
  assign N7 = N161;
  assign N8 = N163;
  assign N9 = N165;
  assign N10 = N174;
  assign N179 = (N0)? 1'b0 : 
                (N1)? 1'b0 : 
                (N2)? 1'b0 : 
                (N3)? 1'b0 : 
                (N4)? 1'b0 : 
                (N5)? 1'b0 : 
                (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b1 : 1'b0;
  assign { N183, N182, N181, N180 } = (N11)? { N178, N177, N176, N175 } : 
                                      (N132)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = N131;
  assign N184 = (N11)? N179 : 
                (N132)? 1'b1 : 1'b0;
  assign { N231, N230, N229 } = (N12)? { 1'b0, 1'b0, 1'b0 } : 
                                (N13)? { 1'b0, 1'b0, 1'b1 } : 
                                (N14)? { 1'b1, 1'b0, 1'b1 } : 
                                (N15)? { 1'b1, 1'b0, 1'b1 } : 
                                (N16)? { 1'b0, 1'b1, 1'b0 } : 
                                (N17)? { 1'b0, 1'b1, 1'b1 } : 
                                (N18)? { 1'b1, 1'b0, 1'b0 } : 
                                (N19)? { 1'b1, 1'b1, 1'b0 } : 
                                (N20)? { 1'b1, 1'b1, 1'b1 } : 
                                (N228)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = N191;
  assign N13 = N196;
  assign N14 = N202;
  assign N15 = N212;
  assign N16 = N213;
  assign N17 = N214;
  assign N18 = N215;
  assign N19 = N217;
  assign N20 = N219;
  assign N232 = (N12)? 1'b0 : 
                (N13)? 1'b0 : 
                (N14)? 1'b0 : 
                (N15)? 1'b0 : 
                (N16)? 1'b0 : 
                (N17)? 1'b0 : 
                (N18)? 1'b0 : 
                (N19)? 1'b0 : 
                (N20)? 1'b0 : 
                (N228)? 1'b1 : 1'b0;
  assign { N236, N235, N234, N233 } = (N21)? { N212, N231, N230, N229 } : 
                                      (N187)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = N186;
  assign N237 = (N21)? N232 : 
                (N187)? 1'b1 : 1'b0;
  assign { N256, N255, N254, N253 } = (N22)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                      (N23)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                      (N24)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N25)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                      (N26)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                      (N27)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                      (N28)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = N243;
  assign N23 = N244;
  assign N24 = N246;
  assign N25 = N247;
  assign N26 = N249;
  assign N27 = N250;
  assign N28 = N252;
  assign N257 = (N22)? 1'b0 : 
                (N23)? 1'b0 : 
                (N24)? 1'b0 : 
                (N25)? 1'b0 : 
                (N26)? 1'b0 : 
                (N27)? 1'b0 : 
                (N28)? 1'b1 : 1'b0;
  assign { N261, N260, N259, N258 } = (N29)? { N256, N255, N254, N253 } : 
                                      (N30)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N29 = N241;
  assign N30 = N240;
  assign N262 = (N29)? N257 : 
                (N30)? 1'b1 : 1'b0;
  assign { N270, N269, N268 } = (N22)? { 1'b0, 1'b0, 1'b0 } : 
                                (N23)? { 1'b0, 1'b0, 1'b1 } : 
                                (N31)? { 1'b0, 1'b1, 1'b0 } : 
                                (N24)? { 1'b1, 1'b0, 1'b0 } : 
                                (N25)? { 1'b1, 1'b0, 1'b1 } : 
                                (N26)? { 1'b1, 1'b1, 1'b0 } : 
                                (N32)? { 1'b0, 1'b1, 1'b1 } : 
                                (N27)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N31 = N266;
  assign N32 = N267;
  assign N271 = (N22)? 1'b0 : 
                (N23)? 1'b0 : 
                (N31)? 1'b0 : 
                (N24)? 1'b0 : 
                (N25)? 1'b0 : 
                (N26)? 1'b0 : 
                (N32)? 1'b0 : 
                (N27)? 1'b1 : 1'b0;
  assign { N274, N273, N272 } = (N33)? { N270, N269, N268 } : 
                                (N34)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N33 = N265;
  assign N34 = N264;
  assign N275 = (N33)? N271 : 
                (N34)? 1'b1 : 1'b0;
  assign { N290, N289 } = (N35)? { 1'b0, 1'b0 } : 
                          (N36)? { 1'b0, 1'b1 } : 
                          (N37)? { 1'b1, 1'b0 } : 
                          (N38)? { 1'b1, 1'b1 } : 1'b0;
  assign N35 = N285;
  assign N36 = N286;
  assign N37 = N287;
  assign N38 = N288;
  assign { N292, N291 } = (N39)? { N290, N289 } : 
                          (N282)? { 1'b0, 1'b0 } : 1'b0;
  assign N39 = N281;
  assign N293 = ~N281;
  assign { N319, N318, N317, N314, N313, N312, N311, N310, N309, N308 } = (N40)? { 1'b1, 1'b0, 1'b1, N350, N183, N182, N181, N180, 1'b0, 1'b0 } : 
                                                                          (N41)? { 1'b1, 1'b0, 1'b1, N357, N236, N235, N234, N233, 1'b1, 1'b0 } : 
                                                                          (N42)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                                          (N43)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                                          (N44)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                                          (N45)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                                          (N46)? { 1'b1, 1'b0, 1'b0, 1'b0, N261, N260, N259, N258, 1'b0, 1'b0 } : 
                                                                          (N47)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, N274, N273, N272, 1'b0, 1'b0 } : 
                                                                          (N48)? { 1'b0, 1'b1, 1'b0, 1'b0, N281, 1'b0, N292, N291, 1'b0, 1'b0 } : 
                                                                          (N49)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N50)? { 1'b1, 1'b0, N307, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N51)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = N63;
  assign N41 = N69;
  assign N42 = N71;
  assign N43 = N73;
  assign N44 = N78;
  assign N45 = N82;
  assign N46 = N84;
  assign N47 = N90;
  assign N48 = N93;
  assign N49 = N96;
  assign N50 = N99;
  assign N51 = N116;
  assign N316 = (N50)? N307 : 
                (N315)? 1'b0 : 1'b0;
  assign N320 = (N40)? N184 : 
                (N41)? N237 : 
                (N42)? 1'b0 : 
                (N43)? 1'b0 : 
                (N44)? 1'b0 : 
                (N45)? 1'b0 : 
                (N46)? N262 : 
                (N47)? N275 : 
                (N48)? N293 : 
                (N49)? 1'b0 : 
                (N50)? N306 : 
                (N51)? 1'b1 : 1'b0;
  assign { N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321 } = (N52)? { N319, N318, N317, N316, N93, N90, N84, N314, N313, N312, N311, N310, N73, N309, N82, N308 } : 
                                                                                                              (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N52 = N54;
  assign illegal_instr_o = (N52)? N320 : 
                           (N55)? 1'b1 : 1'b0;
  assign decode_o[42] = ~decode_o[38];
  assign { decode_o[41:39], decode_o[37:37], decode_o[35:35], decode_o[33:33], decode_o[31:29], decode_o[25:0] } = (N53)? { fe_nop_v_i, be_nop_v_i, me_nop_v_i, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                   (N338)? { 1'b0, 1'b0, 1'b0, N336, N335, N334, N333, N332, N331, N321, N330, N329, N328, N327, N326, N325, instr_i[19:15], instr_i[24:20], instr_i[11:7], N324, N323, N322, N321 } : 1'b0;
  assign N53 = decode_o[38];
  assign N55 = ~N54;
  assign N63 = N358 | N359;
  assign N358 = ~N59;
  assign N359 = ~N62;
  assign N69 = N360 | N361;
  assign N360 = ~N66;
  assign N361 = ~N68;
  assign N71 = ~N70;
  assign N73 = ~N72;
  assign N78 = ~N77;
  assign N82 = ~N81;
  assign N84 = ~N83;
  assign N85 = ~instr_i[6];
  assign N86 = ~instr_i[2];
  assign N93 = ~N92;
  assign N96 = ~N95;
  assign N99 = ~N98;
  assign N116 = N101 | N367;
  assign N367 = N102 | N366;
  assign N366 = N104 | N365;
  assign N365 = N107 | N364;
  assign N364 = N110 | N363;
  assign N363 = N112 | N362;
  assign N362 = N114 | N115;
  assign N117 = ~instr_i[31];
  assign N118 = ~instr_i[29];
  assign N119 = ~instr_i[28];
  assign N120 = ~instr_i[27];
  assign N121 = ~instr_i[26];
  assign N122 = ~instr_i[25];
  assign N132 = ~N131;
  assign N136 = N134 | N135;
  assign N140 = N138 | N139;
  assign N144 = N142 | N143;
  assign N148 = N146 | N147;
  assign N152 = N150 | N151;
  assign N153 = ~instr_i[30];
  assign N174 = N167 | N370;
  assign N370 = N169 | N369;
  assign N369 = N170 | N368;
  assign N368 = N171 | N173;
  assign N187 = ~N186;
  assign N191 = N188 | N190;
  assign N196 = N194 | N195;
  assign N202 = N200 | N201;
  assign N212 = N209 | N211;
  assign N220 = N196 | N191;
  assign N221 = N202 | N220;
  assign N222 = N212 | N221;
  assign N223 = N213 | N222;
  assign N224 = N214 | N223;
  assign N225 = N215 | N224;
  assign N226 = N217 | N225;
  assign N227 = N219 | N226;
  assign N228 = ~N227;
  assign N241 = ~N240;
  assign N251 = ~instr_i[14];
  assign N265 = ~N264;
  assign N282 = ~N281;
  assign N283 = ~instr_i[13];
  assign N284 = ~instr_i[12];
  assign N294 = ~instr_i[24];
  assign N295 = ~instr_i[22];
  assign N307 = ~N306;
  assign N315 = N98;
  assign N337 = N372 | illegal_instr_o;
  assign N372 = N371 | me_nop_v_i;
  assign N371 = fe_nop_v_i | be_nop_v_i;
  assign decode_o[38] = N337;
  assign N338 = ~decode_o[38];

endmodule



module bsg_scan_width_p5_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [4:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__4_ = i[0] | 1'b0;
  assign t_1__3_ = i[1] | i[0];
  assign t_1__2_ = i[2] | i[1];
  assign t_1__1_ = i[3] | i[2];
  assign t_1__0_ = i[4] | i[3];
  assign t_2__4_ = t_1__4_ | 1'b0;
  assign t_2__3_ = t_1__3_ | 1'b0;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__4_ | 1'b0;
  assign o[1] = t_2__3_ | 1'b0;
  assign o[2] = t_2__2_ | 1'b0;
  assign o[3] = t_2__1_ | 1'b0;
  assign o[4] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_width_p5_lo_to_hi_p1
(
  i,
  o
);

  input [4:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire N0,N1,N2,N3;
  wire [4:1] scan_lo;

  bsg_scan_width_p5_or_p1_lo_to_hi_p1
  scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[4] = scan_lo[4] & N0;
  assign N0 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N1;
  assign N1 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N2;
  assign N2 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N3;
  assign N3 = ~o[0];

endmodule



module bsg_mux_one_hot_width_p64_els_p5
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [319:0] data_i;
  input [4:0] sel_one_hot_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191;
  wire [319:0] data_masked;
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[4];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[4];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[4];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[4];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[4];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[4];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[4];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[4];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[4];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[4];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[4];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[4];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[4];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[4];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[4];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[4];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[4];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[4];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[4];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[4];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[4];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[4];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[4];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[4];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[4];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[4];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[4];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[4];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[4];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[4];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[4];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[4];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[4];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[4];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[4];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[4];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[4];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[4];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[4];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[4];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[4];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[4];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[4];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[4];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[4];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[4];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[4];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[4];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[4];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[4];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[4];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[4];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[4];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[4];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[4];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[4];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[4];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[4];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[4];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[4];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[4];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[4];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[4];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[64];
  assign N1 = N0 | data_masked[128];
  assign N0 = data_masked[256] | data_masked[192];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[65];
  assign N4 = N3 | data_masked[129];
  assign N3 = data_masked[257] | data_masked[193];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[66];
  assign N7 = N6 | data_masked[130];
  assign N6 = data_masked[258] | data_masked[194];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[67];
  assign N10 = N9 | data_masked[131];
  assign N9 = data_masked[259] | data_masked[195];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[68];
  assign N13 = N12 | data_masked[132];
  assign N12 = data_masked[260] | data_masked[196];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[69];
  assign N16 = N15 | data_masked[133];
  assign N15 = data_masked[261] | data_masked[197];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[70];
  assign N19 = N18 | data_masked[134];
  assign N18 = data_masked[262] | data_masked[198];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[71];
  assign N22 = N21 | data_masked[135];
  assign N21 = data_masked[263] | data_masked[199];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[72];
  assign N25 = N24 | data_masked[136];
  assign N24 = data_masked[264] | data_masked[200];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[73];
  assign N28 = N27 | data_masked[137];
  assign N27 = data_masked[265] | data_masked[201];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[74];
  assign N31 = N30 | data_masked[138];
  assign N30 = data_masked[266] | data_masked[202];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[75];
  assign N34 = N33 | data_masked[139];
  assign N33 = data_masked[267] | data_masked[203];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[76];
  assign N37 = N36 | data_masked[140];
  assign N36 = data_masked[268] | data_masked[204];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[77];
  assign N40 = N39 | data_masked[141];
  assign N39 = data_masked[269] | data_masked[205];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[78];
  assign N43 = N42 | data_masked[142];
  assign N42 = data_masked[270] | data_masked[206];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[79];
  assign N46 = N45 | data_masked[143];
  assign N45 = data_masked[271] | data_masked[207];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[80];
  assign N49 = N48 | data_masked[144];
  assign N48 = data_masked[272] | data_masked[208];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[81];
  assign N52 = N51 | data_masked[145];
  assign N51 = data_masked[273] | data_masked[209];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[82];
  assign N55 = N54 | data_masked[146];
  assign N54 = data_masked[274] | data_masked[210];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[83];
  assign N58 = N57 | data_masked[147];
  assign N57 = data_masked[275] | data_masked[211];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[84];
  assign N61 = N60 | data_masked[148];
  assign N60 = data_masked[276] | data_masked[212];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[85];
  assign N64 = N63 | data_masked[149];
  assign N63 = data_masked[277] | data_masked[213];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[86];
  assign N67 = N66 | data_masked[150];
  assign N66 = data_masked[278] | data_masked[214];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[87];
  assign N70 = N69 | data_masked[151];
  assign N69 = data_masked[279] | data_masked[215];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[88];
  assign N73 = N72 | data_masked[152];
  assign N72 = data_masked[280] | data_masked[216];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[89];
  assign N76 = N75 | data_masked[153];
  assign N75 = data_masked[281] | data_masked[217];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[90];
  assign N79 = N78 | data_masked[154];
  assign N78 = data_masked[282] | data_masked[218];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[91];
  assign N82 = N81 | data_masked[155];
  assign N81 = data_masked[283] | data_masked[219];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[92];
  assign N85 = N84 | data_masked[156];
  assign N84 = data_masked[284] | data_masked[220];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[93];
  assign N88 = N87 | data_masked[157];
  assign N87 = data_masked[285] | data_masked[221];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[94];
  assign N91 = N90 | data_masked[158];
  assign N90 = data_masked[286] | data_masked[222];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[95];
  assign N94 = N93 | data_masked[159];
  assign N93 = data_masked[287] | data_masked[223];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[96];
  assign N97 = N96 | data_masked[160];
  assign N96 = data_masked[288] | data_masked[224];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[97];
  assign N100 = N99 | data_masked[161];
  assign N99 = data_masked[289] | data_masked[225];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[98];
  assign N103 = N102 | data_masked[162];
  assign N102 = data_masked[290] | data_masked[226];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[99];
  assign N106 = N105 | data_masked[163];
  assign N105 = data_masked[291] | data_masked[227];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[100];
  assign N109 = N108 | data_masked[164];
  assign N108 = data_masked[292] | data_masked[228];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[101];
  assign N112 = N111 | data_masked[165];
  assign N111 = data_masked[293] | data_masked[229];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[102];
  assign N115 = N114 | data_masked[166];
  assign N114 = data_masked[294] | data_masked[230];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[103];
  assign N118 = N117 | data_masked[167];
  assign N117 = data_masked[295] | data_masked[231];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[104];
  assign N121 = N120 | data_masked[168];
  assign N120 = data_masked[296] | data_masked[232];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[105];
  assign N124 = N123 | data_masked[169];
  assign N123 = data_masked[297] | data_masked[233];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[106];
  assign N127 = N126 | data_masked[170];
  assign N126 = data_masked[298] | data_masked[234];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[107];
  assign N130 = N129 | data_masked[171];
  assign N129 = data_masked[299] | data_masked[235];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[108];
  assign N133 = N132 | data_masked[172];
  assign N132 = data_masked[300] | data_masked[236];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[109];
  assign N136 = N135 | data_masked[173];
  assign N135 = data_masked[301] | data_masked[237];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[110];
  assign N139 = N138 | data_masked[174];
  assign N138 = data_masked[302] | data_masked[238];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[111];
  assign N142 = N141 | data_masked[175];
  assign N141 = data_masked[303] | data_masked[239];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[112];
  assign N145 = N144 | data_masked[176];
  assign N144 = data_masked[304] | data_masked[240];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[113];
  assign N148 = N147 | data_masked[177];
  assign N147 = data_masked[305] | data_masked[241];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[114];
  assign N151 = N150 | data_masked[178];
  assign N150 = data_masked[306] | data_masked[242];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[115];
  assign N154 = N153 | data_masked[179];
  assign N153 = data_masked[307] | data_masked[243];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[116];
  assign N157 = N156 | data_masked[180];
  assign N156 = data_masked[308] | data_masked[244];
  assign data_o[53] = N161 | data_masked[53];
  assign N161 = N160 | data_masked[117];
  assign N160 = N159 | data_masked[181];
  assign N159 = data_masked[309] | data_masked[245];
  assign data_o[54] = N164 | data_masked[54];
  assign N164 = N163 | data_masked[118];
  assign N163 = N162 | data_masked[182];
  assign N162 = data_masked[310] | data_masked[246];
  assign data_o[55] = N167 | data_masked[55];
  assign N167 = N166 | data_masked[119];
  assign N166 = N165 | data_masked[183];
  assign N165 = data_masked[311] | data_masked[247];
  assign data_o[56] = N170 | data_masked[56];
  assign N170 = N169 | data_masked[120];
  assign N169 = N168 | data_masked[184];
  assign N168 = data_masked[312] | data_masked[248];
  assign data_o[57] = N173 | data_masked[57];
  assign N173 = N172 | data_masked[121];
  assign N172 = N171 | data_masked[185];
  assign N171 = data_masked[313] | data_masked[249];
  assign data_o[58] = N176 | data_masked[58];
  assign N176 = N175 | data_masked[122];
  assign N175 = N174 | data_masked[186];
  assign N174 = data_masked[314] | data_masked[250];
  assign data_o[59] = N179 | data_masked[59];
  assign N179 = N178 | data_masked[123];
  assign N178 = N177 | data_masked[187];
  assign N177 = data_masked[315] | data_masked[251];
  assign data_o[60] = N182 | data_masked[60];
  assign N182 = N181 | data_masked[124];
  assign N181 = N180 | data_masked[188];
  assign N180 = data_masked[316] | data_masked[252];
  assign data_o[61] = N185 | data_masked[61];
  assign N185 = N184 | data_masked[125];
  assign N184 = N183 | data_masked[189];
  assign N183 = data_masked[317] | data_masked[253];
  assign data_o[62] = N188 | data_masked[62];
  assign N188 = N187 | data_masked[126];
  assign N187 = N186 | data_masked[190];
  assign N186 = data_masked[318] | data_masked[254];
  assign data_o[63] = N191 | data_masked[63];
  assign N191 = N190 | data_masked[127];
  assign N190 = N189 | data_masked[191];
  assign N189 = data_masked[319] | data_masked[255];

endmodule



module bsg_crossbar_o_by_i_i_els_p5_o_els_p1_width_p64
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [319:0] i;
  input [4:0] sel_oi_one_hot_i;
  output [63:0] o;
  wire [63:0] o;

  bsg_mux_one_hot_width_p64_els_p5
  genblk1_0__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i),
    .data_o(o)
  );


endmodule



module bp_be_bypass_fwd_els_p4
(
  id_rs1_v_i,
  id_rs1_addr_i,
  id_rs1_i,
  id_rs2_v_i,
  id_rs2_addr_i,
  id_rs2_i,
  fwd_rd_v_i,
  fwd_rd_addr_i,
  fwd_rd_i,
  bypass_rs1_o,
  bypass_rs2_o
);

  input [4:0] id_rs1_addr_i;
  input [63:0] id_rs1_i;
  input [4:0] id_rs2_addr_i;
  input [63:0] id_rs2_i;
  input [3:0] fwd_rd_v_i;
  input [19:0] fwd_rd_addr_i;
  input [255:0] fwd_rd_i;
  output [63:0] bypass_rs1_o;
  output [63:0] bypass_rs2_o;
  input id_rs1_v_i;
  input id_rs2_v_i;
  wire [63:0] bypass_rs1_o,bypass_rs2_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55;
  wire [3:0] rs1_match_vector,rs2_match_vector;
  wire [4:0] rs1_match_vector_onehot,rs2_match_vector_onehot;

  bsg_priority_encode_one_hot_out_width_p5_lo_to_hi_p1
  bypass_match_one_hot_rs1
  (
    .i({ 1'b1, rs1_match_vector }),
    .o(rs1_match_vector_onehot)
  );


  bsg_priority_encode_one_hot_out_width_p5_lo_to_hi_p1
  bypass_match_one_hot_rs2
  (
    .i({ 1'b1, rs2_match_vector }),
    .o(rs2_match_vector_onehot)
  );


  bsg_crossbar_o_by_i_i_els_p5_o_els_p1_width_p64
  bypass_rs1_crossbar
  (
    .i({ id_rs1_i, fwd_rd_i }),
    .sel_oi_one_hot_i(rs1_match_vector_onehot),
    .o(bypass_rs1_o)
  );


  bsg_crossbar_o_by_i_i_els_p5_o_els_p1_width_p64
  bypass_rs2_crossbar
  (
    .i({ id_rs2_i, fwd_rd_i }),
    .sel_oi_one_hot_i(rs2_match_vector_onehot),
    .o(bypass_rs2_o)
  );

  assign N0 = id_rs1_addr_i == fwd_rd_addr_i[4:0];
  assign N1 = id_rs2_addr_i == fwd_rd_addr_i[4:0];
  assign N2 = id_rs1_addr_i == fwd_rd_addr_i[9:5];
  assign N3 = id_rs2_addr_i == fwd_rd_addr_i[9:5];
  assign N4 = id_rs1_addr_i == fwd_rd_addr_i[14:10];
  assign N5 = id_rs2_addr_i == fwd_rd_addr_i[14:10];
  assign N6 = id_rs1_addr_i == fwd_rd_addr_i[19:15];
  assign N7 = id_rs2_addr_i == fwd_rd_addr_i[19:15];
  assign N8 = id_rs1_addr_i[3] | id_rs1_addr_i[4];
  assign N9 = id_rs1_addr_i[2] | N8;
  assign N10 = id_rs1_addr_i[1] | N9;
  assign N11 = id_rs1_addr_i[0] | N10;
  assign N12 = id_rs1_addr_i[3] | id_rs1_addr_i[4];
  assign N13 = id_rs1_addr_i[2] | N12;
  assign N14 = id_rs1_addr_i[1] | N13;
  assign N15 = id_rs1_addr_i[0] | N14;
  assign N16 = id_rs1_addr_i[3] | id_rs1_addr_i[4];
  assign N17 = id_rs1_addr_i[2] | N16;
  assign N18 = id_rs1_addr_i[1] | N17;
  assign N19 = id_rs1_addr_i[0] | N18;
  assign N20 = id_rs1_addr_i[3] | id_rs1_addr_i[4];
  assign N21 = id_rs1_addr_i[2] | N20;
  assign N22 = id_rs1_addr_i[1] | N21;
  assign N23 = id_rs1_addr_i[0] | N22;
  assign N24 = id_rs2_addr_i[3] | id_rs2_addr_i[4];
  assign N25 = id_rs2_addr_i[2] | N24;
  assign N26 = id_rs2_addr_i[1] | N25;
  assign N27 = id_rs2_addr_i[0] | N26;
  assign N28 = id_rs2_addr_i[3] | id_rs2_addr_i[4];
  assign N29 = id_rs2_addr_i[2] | N28;
  assign N30 = id_rs2_addr_i[1] | N29;
  assign N31 = id_rs2_addr_i[0] | N30;
  assign N32 = id_rs2_addr_i[3] | id_rs2_addr_i[4];
  assign N33 = id_rs2_addr_i[2] | N32;
  assign N34 = id_rs2_addr_i[1] | N33;
  assign N35 = id_rs2_addr_i[0] | N34;
  assign N36 = id_rs2_addr_i[3] | id_rs2_addr_i[4];
  assign N37 = id_rs2_addr_i[2] | N36;
  assign N38 = id_rs2_addr_i[1] | N37;
  assign N39 = id_rs2_addr_i[0] | N38;
  assign rs1_match_vector[0] = N41 & N23;
  assign N41 = N0 & N40;
  assign N40 = id_rs1_v_i & fwd_rd_v_i[0];
  assign rs2_match_vector[0] = N43 & N39;
  assign N43 = N1 & N42;
  assign N42 = id_rs2_v_i & fwd_rd_v_i[0];
  assign rs1_match_vector[1] = N45 & N19;
  assign N45 = N2 & N44;
  assign N44 = id_rs1_v_i & fwd_rd_v_i[1];
  assign rs2_match_vector[1] = N47 & N35;
  assign N47 = N3 & N46;
  assign N46 = id_rs2_v_i & fwd_rd_v_i[1];
  assign rs1_match_vector[2] = N49 & N15;
  assign N49 = N4 & N48;
  assign N48 = id_rs1_v_i & fwd_rd_v_i[2];
  assign rs2_match_vector[2] = N51 & N31;
  assign N51 = N5 & N50;
  assign N50 = id_rs2_v_i & fwd_rd_v_i[2];
  assign rs1_match_vector[3] = N53 & N11;
  assign N53 = N6 & N52;
  assign N52 = id_rs1_v_i & fwd_rd_v_i[3];
  assign rs2_match_vector[3] = N55 & N27;
  assign N55 = N7 & N54;
  assign N54 = id_rs2_v_i & fwd_rd_v_i[3];

endmodule



module bp_be_int_alu
(
  src1_i,
  src2_i,
  op_i,
  opw_v_i,
  result_o
);

  input [63:0] src1_i;
  input [63:0] src2_i;
  input [3:0] op_i;
  output [63:0] result_o;
  input opw_v_i;
  wire [63:0] result_o,result_sgn;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795;
  wire [31:0] resultw_sgn;
  assign N27 = N231 & N35;
  assign N28 = N272 | op_i[0];
  assign N30 = N248 | N35;
  assign N32 = N237 | N35;
  assign N34 = N256 & op_i[0];
  assign N36 = N272 | N35;
  assign N37 = op_i[2] & N35;
  assign { N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103 } = src1_i[31:0] << src2_i[4:0];
  assign { N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135 } = src1_i[31:0] >> src2_i[4:0];
  assign { N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167 } = $signed(src1_i[31:0]) >>> src2_i[4:0];
  assign N231 = N271 & N236;
  assign N232 = N241 & N35;
  assign N233 = N231 & N232;
  assign N234 = N272 | N238;
  assign N237 = op_i[3] | N236;
  assign N238 = op_i[1] | op_i[0];
  assign N239 = N237 | N238;
  assign N242 = N241 | op_i[0];
  assign N243 = N237 | N242;
  assign N245 = N241 | N35;
  assign N246 = N237 | N245;
  assign N248 = op_i[3] | op_i[2];
  assign N249 = N248 | N273;
  assign N251 = N237 | N273;
  assign N253 = N271 | N236;
  assign N254 = N253 | N273;
  assign N256 = op_i[3] & op_i[2];
  assign N257 = op_i[1] & op_i[0];
  assign N258 = N256 & N257;
  assign N259 = N248 | N242;
  assign N261 = N272 | N242;
  assign N263 = N253 | N238;
  assign N265 = N253 | N242;
  assign N267 = N248 | N245;
  assign N269 = N272 | N245;
  assign N272 = N271 | op_i[2];
  assign N273 = op_i[1] | N35;
  assign N274 = N272 | N273;
  assign { N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596 } = src1_i << src2_i[5:0];
  assign { N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660 } = src1_i >> src2_i[5:0];
  assign { N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724 } = $signed(src1_i) >>> src2_i[5:0];
  assign N788 = $signed(src1_i) < $signed(src2_i);
  assign N789 = $signed(src1_i) >= $signed(src2_i);
  assign N790 = src1_i == src2_i;
  assign N791 = src1_i != src2_i;
  assign N792 = src1_i < src2_i;
  assign N793 = src1_i >= src2_i;
  assign { N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276 } = $signed(src1_i) + $signed(src2_i);
  assign { N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39 } = $signed(src1_i[31:0]) + $signed(src2_i[31:0]);
  assign { N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340 } = $signed(src1_i) - $signed(src2_i);
  assign { N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71 } = $signed(src1_i[31:0]) - $signed(src2_i[31:0]);
  assign { N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199 } = (N0)? { N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39 } : 
                                                                                                                                                                                                              (N1)? { N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71 } : 
                                                                                                                                                                                                              (N2)? { N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103 } : 
                                                                                                                                                                                                              (N3)? { N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135 } : 
                                                                                                                                                                                                              (N4)? { N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167 } : 
                                                                                                                                                                                                              (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N27;
  assign N1 = N29;
  assign N2 = N31;
  assign N3 = N33;
  assign N4 = N34;
  assign N5 = N38;
  assign resultw_sgn = (N6)? { N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199 } : 
                       (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = N241;
  assign N7 = op_i[1];
  assign result_sgn = (N8)? { N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276 } : 
                      (N9)? { N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340 } : 
                      (N10)? { N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467 } : 
                      (N11)? { N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531 } : 
                      (N12)? { N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595 } : 
                      (N13)? { N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596 } : 
                      (N14)? { N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660 } : 
                      (N15)? { N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724 } : 
                      (N16)? src2_i : 
                      (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N788 } : 
                      (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N789 } : 
                      (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N790 } : 
                      (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N791 } : 
                      (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N792 } : 
                      (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N793 } : 
                      (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N233;
  assign N9 = N235;
  assign N10 = N240;
  assign N11 = N244;
  assign N12 = N247;
  assign N13 = N250;
  assign N14 = N252;
  assign N15 = N255;
  assign N16 = N258;
  assign N17 = N260;
  assign N18 = N262;
  assign N19 = N264;
  assign N20 = N266;
  assign N21 = N268;
  assign N22 = N270;
  assign N23 = N275;
  assign result_o = (N24)? { resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn } : 
                    (N25)? result_sgn : 1'b0;
  assign N24 = opw_v_i;
  assign N25 = N794;
  assign N26 = N241;
  assign N29 = ~N28;
  assign N31 = ~N30;
  assign N33 = ~N32;
  assign N35 = ~op_i[0];
  assign N38 = N795 | N37;
  assign N795 = ~N36;
  assign N235 = ~N234;
  assign N236 = ~op_i[2];
  assign N240 = ~N239;
  assign N241 = ~op_i[1];
  assign N244 = ~N243;
  assign N247 = ~N246;
  assign N250 = ~N249;
  assign N252 = ~N251;
  assign N255 = ~N254;
  assign N260 = ~N259;
  assign N262 = ~N261;
  assign N264 = ~N263;
  assign N266 = ~N265;
  assign N268 = ~N267;
  assign N270 = ~N269;
  assign N271 = ~op_i[3];
  assign N275 = ~N274;
  assign N404 = src1_i[63] ^ src2_i[63];
  assign N405 = src1_i[62] ^ src2_i[62];
  assign N406 = src1_i[61] ^ src2_i[61];
  assign N407 = src1_i[60] ^ src2_i[60];
  assign N408 = src1_i[59] ^ src2_i[59];
  assign N409 = src1_i[58] ^ src2_i[58];
  assign N410 = src1_i[57] ^ src2_i[57];
  assign N411 = src1_i[56] ^ src2_i[56];
  assign N412 = src1_i[55] ^ src2_i[55];
  assign N413 = src1_i[54] ^ src2_i[54];
  assign N414 = src1_i[53] ^ src2_i[53];
  assign N415 = src1_i[52] ^ src2_i[52];
  assign N416 = src1_i[51] ^ src2_i[51];
  assign N417 = src1_i[50] ^ src2_i[50];
  assign N418 = src1_i[49] ^ src2_i[49];
  assign N419 = src1_i[48] ^ src2_i[48];
  assign N420 = src1_i[47] ^ src2_i[47];
  assign N421 = src1_i[46] ^ src2_i[46];
  assign N422 = src1_i[45] ^ src2_i[45];
  assign N423 = src1_i[44] ^ src2_i[44];
  assign N424 = src1_i[43] ^ src2_i[43];
  assign N425 = src1_i[42] ^ src2_i[42];
  assign N426 = src1_i[41] ^ src2_i[41];
  assign N427 = src1_i[40] ^ src2_i[40];
  assign N428 = src1_i[39] ^ src2_i[39];
  assign N429 = src1_i[38] ^ src2_i[38];
  assign N430 = src1_i[37] ^ src2_i[37];
  assign N431 = src1_i[36] ^ src2_i[36];
  assign N432 = src1_i[35] ^ src2_i[35];
  assign N433 = src1_i[34] ^ src2_i[34];
  assign N434 = src1_i[33] ^ src2_i[33];
  assign N435 = src1_i[32] ^ src2_i[32];
  assign N436 = src1_i[31] ^ src2_i[31];
  assign N437 = src1_i[30] ^ src2_i[30];
  assign N438 = src1_i[29] ^ src2_i[29];
  assign N439 = src1_i[28] ^ src2_i[28];
  assign N440 = src1_i[27] ^ src2_i[27];
  assign N441 = src1_i[26] ^ src2_i[26];
  assign N442 = src1_i[25] ^ src2_i[25];
  assign N443 = src1_i[24] ^ src2_i[24];
  assign N444 = src1_i[23] ^ src2_i[23];
  assign N445 = src1_i[22] ^ src2_i[22];
  assign N446 = src1_i[21] ^ src2_i[21];
  assign N447 = src1_i[20] ^ src2_i[20];
  assign N448 = src1_i[19] ^ src2_i[19];
  assign N449 = src1_i[18] ^ src2_i[18];
  assign N450 = src1_i[17] ^ src2_i[17];
  assign N451 = src1_i[16] ^ src2_i[16];
  assign N452 = src1_i[15] ^ src2_i[15];
  assign N453 = src1_i[14] ^ src2_i[14];
  assign N454 = src1_i[13] ^ src2_i[13];
  assign N455 = src1_i[12] ^ src2_i[12];
  assign N456 = src1_i[11] ^ src2_i[11];
  assign N457 = src1_i[10] ^ src2_i[10];
  assign N458 = src1_i[9] ^ src2_i[9];
  assign N459 = src1_i[8] ^ src2_i[8];
  assign N460 = src1_i[7] ^ src2_i[7];
  assign N461 = src1_i[6] ^ src2_i[6];
  assign N462 = src1_i[5] ^ src2_i[5];
  assign N463 = src1_i[4] ^ src2_i[4];
  assign N464 = src1_i[3] ^ src2_i[3];
  assign N465 = src1_i[2] ^ src2_i[2];
  assign N466 = src1_i[1] ^ src2_i[1];
  assign N467 = src1_i[0] ^ src2_i[0];
  assign N468 = src1_i[63] | src2_i[63];
  assign N469 = src1_i[62] | src2_i[62];
  assign N470 = src1_i[61] | src2_i[61];
  assign N471 = src1_i[60] | src2_i[60];
  assign N472 = src1_i[59] | src2_i[59];
  assign N473 = src1_i[58] | src2_i[58];
  assign N474 = src1_i[57] | src2_i[57];
  assign N475 = src1_i[56] | src2_i[56];
  assign N476 = src1_i[55] | src2_i[55];
  assign N477 = src1_i[54] | src2_i[54];
  assign N478 = src1_i[53] | src2_i[53];
  assign N479 = src1_i[52] | src2_i[52];
  assign N480 = src1_i[51] | src2_i[51];
  assign N481 = src1_i[50] | src2_i[50];
  assign N482 = src1_i[49] | src2_i[49];
  assign N483 = src1_i[48] | src2_i[48];
  assign N484 = src1_i[47] | src2_i[47];
  assign N485 = src1_i[46] | src2_i[46];
  assign N486 = src1_i[45] | src2_i[45];
  assign N487 = src1_i[44] | src2_i[44];
  assign N488 = src1_i[43] | src2_i[43];
  assign N489 = src1_i[42] | src2_i[42];
  assign N490 = src1_i[41] | src2_i[41];
  assign N491 = src1_i[40] | src2_i[40];
  assign N492 = src1_i[39] | src2_i[39];
  assign N493 = src1_i[38] | src2_i[38];
  assign N494 = src1_i[37] | src2_i[37];
  assign N495 = src1_i[36] | src2_i[36];
  assign N496 = src1_i[35] | src2_i[35];
  assign N497 = src1_i[34] | src2_i[34];
  assign N498 = src1_i[33] | src2_i[33];
  assign N499 = src1_i[32] | src2_i[32];
  assign N500 = src1_i[31] | src2_i[31];
  assign N501 = src1_i[30] | src2_i[30];
  assign N502 = src1_i[29] | src2_i[29];
  assign N503 = src1_i[28] | src2_i[28];
  assign N504 = src1_i[27] | src2_i[27];
  assign N505 = src1_i[26] | src2_i[26];
  assign N506 = src1_i[25] | src2_i[25];
  assign N507 = src1_i[24] | src2_i[24];
  assign N508 = src1_i[23] | src2_i[23];
  assign N509 = src1_i[22] | src2_i[22];
  assign N510 = src1_i[21] | src2_i[21];
  assign N511 = src1_i[20] | src2_i[20];
  assign N512 = src1_i[19] | src2_i[19];
  assign N513 = src1_i[18] | src2_i[18];
  assign N514 = src1_i[17] | src2_i[17];
  assign N515 = src1_i[16] | src2_i[16];
  assign N516 = src1_i[15] | src2_i[15];
  assign N517 = src1_i[14] | src2_i[14];
  assign N518 = src1_i[13] | src2_i[13];
  assign N519 = src1_i[12] | src2_i[12];
  assign N520 = src1_i[11] | src2_i[11];
  assign N521 = src1_i[10] | src2_i[10];
  assign N522 = src1_i[9] | src2_i[9];
  assign N523 = src1_i[8] | src2_i[8];
  assign N524 = src1_i[7] | src2_i[7];
  assign N525 = src1_i[6] | src2_i[6];
  assign N526 = src1_i[5] | src2_i[5];
  assign N527 = src1_i[4] | src2_i[4];
  assign N528 = src1_i[3] | src2_i[3];
  assign N529 = src1_i[2] | src2_i[2];
  assign N530 = src1_i[1] | src2_i[1];
  assign N531 = src1_i[0] | src2_i[0];
  assign N532 = src1_i[63] & src2_i[63];
  assign N533 = src1_i[62] & src2_i[62];
  assign N534 = src1_i[61] & src2_i[61];
  assign N535 = src1_i[60] & src2_i[60];
  assign N536 = src1_i[59] & src2_i[59];
  assign N537 = src1_i[58] & src2_i[58];
  assign N538 = src1_i[57] & src2_i[57];
  assign N539 = src1_i[56] & src2_i[56];
  assign N540 = src1_i[55] & src2_i[55];
  assign N541 = src1_i[54] & src2_i[54];
  assign N542 = src1_i[53] & src2_i[53];
  assign N543 = src1_i[52] & src2_i[52];
  assign N544 = src1_i[51] & src2_i[51];
  assign N545 = src1_i[50] & src2_i[50];
  assign N546 = src1_i[49] & src2_i[49];
  assign N547 = src1_i[48] & src2_i[48];
  assign N548 = src1_i[47] & src2_i[47];
  assign N549 = src1_i[46] & src2_i[46];
  assign N550 = src1_i[45] & src2_i[45];
  assign N551 = src1_i[44] & src2_i[44];
  assign N552 = src1_i[43] & src2_i[43];
  assign N553 = src1_i[42] & src2_i[42];
  assign N554 = src1_i[41] & src2_i[41];
  assign N555 = src1_i[40] & src2_i[40];
  assign N556 = src1_i[39] & src2_i[39];
  assign N557 = src1_i[38] & src2_i[38];
  assign N558 = src1_i[37] & src2_i[37];
  assign N559 = src1_i[36] & src2_i[36];
  assign N560 = src1_i[35] & src2_i[35];
  assign N561 = src1_i[34] & src2_i[34];
  assign N562 = src1_i[33] & src2_i[33];
  assign N563 = src1_i[32] & src2_i[32];
  assign N564 = src1_i[31] & src2_i[31];
  assign N565 = src1_i[30] & src2_i[30];
  assign N566 = src1_i[29] & src2_i[29];
  assign N567 = src1_i[28] & src2_i[28];
  assign N568 = src1_i[27] & src2_i[27];
  assign N569 = src1_i[26] & src2_i[26];
  assign N570 = src1_i[25] & src2_i[25];
  assign N571 = src1_i[24] & src2_i[24];
  assign N572 = src1_i[23] & src2_i[23];
  assign N573 = src1_i[22] & src2_i[22];
  assign N574 = src1_i[21] & src2_i[21];
  assign N575 = src1_i[20] & src2_i[20];
  assign N576 = src1_i[19] & src2_i[19];
  assign N577 = src1_i[18] & src2_i[18];
  assign N578 = src1_i[17] & src2_i[17];
  assign N579 = src1_i[16] & src2_i[16];
  assign N580 = src1_i[15] & src2_i[15];
  assign N581 = src1_i[14] & src2_i[14];
  assign N582 = src1_i[13] & src2_i[13];
  assign N583 = src1_i[12] & src2_i[12];
  assign N584 = src1_i[11] & src2_i[11];
  assign N585 = src1_i[10] & src2_i[10];
  assign N586 = src1_i[9] & src2_i[9];
  assign N587 = src1_i[8] & src2_i[8];
  assign N588 = src1_i[7] & src2_i[7];
  assign N589 = src1_i[6] & src2_i[6];
  assign N590 = src1_i[5] & src2_i[5];
  assign N591 = src1_i[4] & src2_i[4];
  assign N592 = src1_i[3] & src2_i[3];
  assign N593 = src1_i[2] & src2_i[2];
  assign N594 = src1_i[1] & src2_i[1];
  assign N595 = src1_i[0] & src2_i[0];
  assign N794 = ~opw_v_i;

endmodule



module bp_be_pipe_int_core_els_p1
(
  clk_i,
  reset_i,
  decode_i,
  pc_i,
  rs1_i,
  rs2_i,
  imm_i,
  exc_i,
  mhartid_i,
  result_o,
  br_tgt_o
);

  input [42:0] decode_i;
  input [63:0] pc_i;
  input [63:0] rs1_i;
  input [63:0] rs2_i;
  input [63:0] imm_i;
  input [6:0] exc_i;
  input [0:0] mhartid_i;
  output [63:0] result_o;
  output [63:0] br_tgt_o;
  input clk_i;
  input reset_i;
  wire [63:0] result_o,br_tgt_o,src1,src2,alu_result,baddr,pc_plus4;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

  bp_be_int_alu
  alu
  (
    .src1_i(src1),
    .src2_i(src2),
    .op_i(decode_i[22:19]),
    .opw_v_i(decode_i[23]),
    .result_o(alu_result)
  );

  assign pc_plus4 = pc_i + { 1'b1, 1'b0, 1'b0 };
  assign br_tgt_o = baddr + imm_i;
  assign src1 = (N0)? pc_i : 
                (N4)? rs1_i : 1'b0;
  assign N0 = decode_i[3];
  assign src2 = (N1)? imm_i : 
                (N5)? rs2_i : 1'b0;
  assign N1 = decode_i[2];
  assign baddr = (N2)? src1 : 
                 (N6)? pc_i : 1'b0;
  assign N2 = decode_i[1];
  assign result_o = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mhartid_i[0:0] } : 
                    (N10)? pc_plus4 : 
                    (N8)? alu_result : 1'b0;
  assign N3 = decode_i[31];
  assign N4 = ~decode_i[3];
  assign N5 = ~decode_i[2];
  assign N6 = ~decode_i[1];
  assign N7 = decode_i[0] | decode_i[31];
  assign N8 = ~N7;
  assign N9 = ~decode_i[31];
  assign N10 = decode_i[0] & N9;

endmodule



module bp_be_pipe_mul
(
  clk_i,
  reset_i,
  decode_i,
  rs1_i,
  rs2_i,
  exc_i,
  result_o
);

  input [42:0] decode_i;
  input [63:0] rs1_i;
  input [63:0] rs2_i;
  input [6:0] exc_i;
  output [63:0] result_o;
  input clk_i;
  input reset_i;
  wire [63:0] result_o;
  assign result_o[0] = 1'b0;
  assign result_o[1] = 1'b0;
  assign result_o[2] = 1'b0;
  assign result_o[3] = 1'b0;
  assign result_o[4] = 1'b0;
  assign result_o[5] = 1'b0;
  assign result_o[6] = 1'b0;
  assign result_o[7] = 1'b0;
  assign result_o[8] = 1'b0;
  assign result_o[9] = 1'b0;
  assign result_o[10] = 1'b0;
  assign result_o[11] = 1'b0;
  assign result_o[12] = 1'b0;
  assign result_o[13] = 1'b0;
  assign result_o[14] = 1'b0;
  assign result_o[15] = 1'b0;
  assign result_o[16] = 1'b0;
  assign result_o[17] = 1'b0;
  assign result_o[18] = 1'b0;
  assign result_o[19] = 1'b0;
  assign result_o[20] = 1'b0;
  assign result_o[21] = 1'b0;
  assign result_o[22] = 1'b0;
  assign result_o[23] = 1'b0;
  assign result_o[24] = 1'b0;
  assign result_o[25] = 1'b0;
  assign result_o[26] = 1'b0;
  assign result_o[27] = 1'b0;
  assign result_o[28] = 1'b0;
  assign result_o[29] = 1'b0;
  assign result_o[30] = 1'b0;
  assign result_o[31] = 1'b0;
  assign result_o[32] = 1'b0;
  assign result_o[33] = 1'b0;
  assign result_o[34] = 1'b0;
  assign result_o[35] = 1'b0;
  assign result_o[36] = 1'b0;
  assign result_o[37] = 1'b0;
  assign result_o[38] = 1'b0;
  assign result_o[39] = 1'b0;
  assign result_o[40] = 1'b0;
  assign result_o[41] = 1'b0;
  assign result_o[42] = 1'b0;
  assign result_o[43] = 1'b0;
  assign result_o[44] = 1'b0;
  assign result_o[45] = 1'b0;
  assign result_o[46] = 1'b0;
  assign result_o[47] = 1'b0;
  assign result_o[48] = 1'b0;
  assign result_o[49] = 1'b0;
  assign result_o[50] = 1'b0;
  assign result_o[51] = 1'b0;
  assign result_o[52] = 1'b0;
  assign result_o[53] = 1'b0;
  assign result_o[54] = 1'b0;
  assign result_o[55] = 1'b0;
  assign result_o[56] = 1'b0;
  assign result_o[57] = 1'b0;
  assign result_o[58] = 1'b0;
  assign result_o[59] = 1'b0;
  assign result_o[60] = 1'b0;
  assign result_o[61] = 1'b0;
  assign result_o[62] = 1'b0;
  assign result_o[63] = 1'b0;

endmodule



module bp_be_pipe_mem_vaddr_width_p56_lce_sets_p64_cce_block_size_in_bytes_p64
(
  clk_i,
  reset_i,
  decode_i,
  rs1_i,
  rs2_i,
  imm_i,
  exc_i,
  mmu_cmd_o,
  mmu_cmd_v_o,
  mmu_cmd_ready_i,
  mmu_resp_i,
  mmu_resp_v_i,
  mmu_resp_ready_o,
  result_o,
  cache_miss_o
);

  input [42:0] decode_i;
  input [63:0] rs1_i;
  input [63:0] rs2_i;
  input [63:0] imm_i;
  input [6:0] exc_i;
  output [123:0] mmu_cmd_o;
  input [70:0] mmu_resp_i;
  output [63:0] result_o;
  input clk_i;
  input reset_i;
  input mmu_cmd_ready_i;
  input mmu_resp_v_i;
  output mmu_cmd_v_o;
  output mmu_resp_ready_o;
  output cache_miss_o;
  wire [123:0] mmu_cmd_o;
  wire [63:0] result_o;
  wire mmu_cmd_v_o,mmu_resp_ready_o,cache_miss_o,N0,N1,N2,N3,N4,N5,N6,N7;
  assign mmu_resp_ready_o = 1'b1;
  assign mmu_cmd_o[123] = decode_i[22];
  assign mmu_cmd_o[122] = decode_i[21];
  assign mmu_cmd_o[121] = decode_i[20];
  assign mmu_cmd_o[120] = decode_i[19];
  assign mmu_cmd_o[63] = rs2_i[63];
  assign mmu_cmd_o[62] = rs2_i[62];
  assign mmu_cmd_o[61] = rs2_i[61];
  assign mmu_cmd_o[60] = rs2_i[60];
  assign mmu_cmd_o[59] = rs2_i[59];
  assign mmu_cmd_o[58] = rs2_i[58];
  assign mmu_cmd_o[57] = rs2_i[57];
  assign mmu_cmd_o[56] = rs2_i[56];
  assign mmu_cmd_o[55] = rs2_i[55];
  assign mmu_cmd_o[54] = rs2_i[54];
  assign mmu_cmd_o[53] = rs2_i[53];
  assign mmu_cmd_o[52] = rs2_i[52];
  assign mmu_cmd_o[51] = rs2_i[51];
  assign mmu_cmd_o[50] = rs2_i[50];
  assign mmu_cmd_o[49] = rs2_i[49];
  assign mmu_cmd_o[48] = rs2_i[48];
  assign mmu_cmd_o[47] = rs2_i[47];
  assign mmu_cmd_o[46] = rs2_i[46];
  assign mmu_cmd_o[45] = rs2_i[45];
  assign mmu_cmd_o[44] = rs2_i[44];
  assign mmu_cmd_o[43] = rs2_i[43];
  assign mmu_cmd_o[42] = rs2_i[42];
  assign mmu_cmd_o[41] = rs2_i[41];
  assign mmu_cmd_o[40] = rs2_i[40];
  assign mmu_cmd_o[39] = rs2_i[39];
  assign mmu_cmd_o[38] = rs2_i[38];
  assign mmu_cmd_o[37] = rs2_i[37];
  assign mmu_cmd_o[36] = rs2_i[36];
  assign mmu_cmd_o[35] = rs2_i[35];
  assign mmu_cmd_o[34] = rs2_i[34];
  assign mmu_cmd_o[33] = rs2_i[33];
  assign mmu_cmd_o[32] = rs2_i[32];
  assign mmu_cmd_o[31] = rs2_i[31];
  assign mmu_cmd_o[30] = rs2_i[30];
  assign mmu_cmd_o[29] = rs2_i[29];
  assign mmu_cmd_o[28] = rs2_i[28];
  assign mmu_cmd_o[27] = rs2_i[27];
  assign mmu_cmd_o[26] = rs2_i[26];
  assign mmu_cmd_o[25] = rs2_i[25];
  assign mmu_cmd_o[24] = rs2_i[24];
  assign mmu_cmd_o[23] = rs2_i[23];
  assign mmu_cmd_o[22] = rs2_i[22];
  assign mmu_cmd_o[21] = rs2_i[21];
  assign mmu_cmd_o[20] = rs2_i[20];
  assign mmu_cmd_o[19] = rs2_i[19];
  assign mmu_cmd_o[18] = rs2_i[18];
  assign mmu_cmd_o[17] = rs2_i[17];
  assign mmu_cmd_o[16] = rs2_i[16];
  assign mmu_cmd_o[15] = rs2_i[15];
  assign mmu_cmd_o[14] = rs2_i[14];
  assign mmu_cmd_o[13] = rs2_i[13];
  assign mmu_cmd_o[12] = rs2_i[12];
  assign mmu_cmd_o[11] = rs2_i[11];
  assign mmu_cmd_o[10] = rs2_i[10];
  assign mmu_cmd_o[9] = rs2_i[9];
  assign mmu_cmd_o[8] = rs2_i[8];
  assign mmu_cmd_o[7] = rs2_i[7];
  assign mmu_cmd_o[6] = rs2_i[6];
  assign mmu_cmd_o[5] = rs2_i[5];
  assign mmu_cmd_o[4] = rs2_i[4];
  assign mmu_cmd_o[3] = rs2_i[3];
  assign mmu_cmd_o[2] = rs2_i[2];
  assign mmu_cmd_o[1] = rs2_i[1];
  assign mmu_cmd_o[0] = rs2_i[0];
  assign result_o[63] = mmu_resp_i[70];
  assign result_o[62] = mmu_resp_i[69];
  assign result_o[61] = mmu_resp_i[68];
  assign result_o[60] = mmu_resp_i[67];
  assign result_o[59] = mmu_resp_i[66];
  assign result_o[58] = mmu_resp_i[65];
  assign result_o[57] = mmu_resp_i[64];
  assign result_o[56] = mmu_resp_i[63];
  assign result_o[55] = mmu_resp_i[62];
  assign result_o[54] = mmu_resp_i[61];
  assign result_o[53] = mmu_resp_i[60];
  assign result_o[52] = mmu_resp_i[59];
  assign result_o[51] = mmu_resp_i[58];
  assign result_o[50] = mmu_resp_i[57];
  assign result_o[49] = mmu_resp_i[56];
  assign result_o[48] = mmu_resp_i[55];
  assign result_o[47] = mmu_resp_i[54];
  assign result_o[46] = mmu_resp_i[53];
  assign result_o[45] = mmu_resp_i[52];
  assign result_o[44] = mmu_resp_i[51];
  assign result_o[43] = mmu_resp_i[50];
  assign result_o[42] = mmu_resp_i[49];
  assign result_o[41] = mmu_resp_i[48];
  assign result_o[40] = mmu_resp_i[47];
  assign result_o[39] = mmu_resp_i[46];
  assign result_o[38] = mmu_resp_i[45];
  assign result_o[37] = mmu_resp_i[44];
  assign result_o[36] = mmu_resp_i[43];
  assign result_o[35] = mmu_resp_i[42];
  assign result_o[34] = mmu_resp_i[41];
  assign result_o[33] = mmu_resp_i[40];
  assign result_o[32] = mmu_resp_i[39];
  assign result_o[31] = mmu_resp_i[38];
  assign result_o[30] = mmu_resp_i[37];
  assign result_o[29] = mmu_resp_i[36];
  assign result_o[28] = mmu_resp_i[35];
  assign result_o[27] = mmu_resp_i[34];
  assign result_o[26] = mmu_resp_i[33];
  assign result_o[25] = mmu_resp_i[32];
  assign result_o[24] = mmu_resp_i[31];
  assign result_o[23] = mmu_resp_i[30];
  assign result_o[22] = mmu_resp_i[29];
  assign result_o[21] = mmu_resp_i[28];
  assign result_o[20] = mmu_resp_i[27];
  assign result_o[19] = mmu_resp_i[26];
  assign result_o[18] = mmu_resp_i[25];
  assign result_o[17] = mmu_resp_i[24];
  assign result_o[16] = mmu_resp_i[23];
  assign result_o[15] = mmu_resp_i[22];
  assign result_o[14] = mmu_resp_i[21];
  assign result_o[13] = mmu_resp_i[20];
  assign result_o[12] = mmu_resp_i[19];
  assign result_o[11] = mmu_resp_i[18];
  assign result_o[10] = mmu_resp_i[17];
  assign result_o[9] = mmu_resp_i[16];
  assign result_o[8] = mmu_resp_i[15];
  assign result_o[7] = mmu_resp_i[14];
  assign result_o[6] = mmu_resp_i[13];
  assign result_o[5] = mmu_resp_i[12];
  assign result_o[4] = mmu_resp_i[11];
  assign result_o[3] = mmu_resp_i[10];
  assign result_o[2] = mmu_resp_i[9];
  assign result_o[1] = mmu_resp_i[8];
  assign result_o[0] = mmu_resp_i[7];
  assign cache_miss_o = mmu_resp_i[0];
  assign mmu_cmd_o[119:64] = rs1_i[55:0] + imm_i[55:0];
  assign mmu_cmd_v_o = N0 & N7;
  assign N0 = decode_i[29] | decode_i[30];
  assign N7 = ~N6;
  assign N6 = N5 | exc_i[0];
  assign N5 = N4 | exc_i[1];
  assign N4 = N3 | exc_i[2];
  assign N3 = N2 | exc_i[3];
  assign N2 = N1 | exc_i[4];
  assign N1 = exc_i[6] | exc_i[5];

endmodule



module bp_be_pipe_fp
(
  clk_i,
  reset_i,
  decode_i,
  rs1_i,
  rs2_i,
  exc_i,
  result_o
);

  input [42:0] decode_i;
  input [63:0] rs1_i;
  input [63:0] rs2_i;
  input [6:0] exc_i;
  output [63:0] result_o;
  input clk_i;
  input reset_i;
  wire [63:0] result_o;
  assign result_o[0] = 1'b0;
  assign result_o[1] = 1'b0;
  assign result_o[2] = 1'b0;
  assign result_o[3] = 1'b0;
  assign result_o[4] = 1'b0;
  assign result_o[5] = 1'b0;
  assign result_o[6] = 1'b0;
  assign result_o[7] = 1'b0;
  assign result_o[8] = 1'b0;
  assign result_o[9] = 1'b0;
  assign result_o[10] = 1'b0;
  assign result_o[11] = 1'b0;
  assign result_o[12] = 1'b0;
  assign result_o[13] = 1'b0;
  assign result_o[14] = 1'b0;
  assign result_o[15] = 1'b0;
  assign result_o[16] = 1'b0;
  assign result_o[17] = 1'b0;
  assign result_o[18] = 1'b0;
  assign result_o[19] = 1'b0;
  assign result_o[20] = 1'b0;
  assign result_o[21] = 1'b0;
  assign result_o[22] = 1'b0;
  assign result_o[23] = 1'b0;
  assign result_o[24] = 1'b0;
  assign result_o[25] = 1'b0;
  assign result_o[26] = 1'b0;
  assign result_o[27] = 1'b0;
  assign result_o[28] = 1'b0;
  assign result_o[29] = 1'b0;
  assign result_o[30] = 1'b0;
  assign result_o[31] = 1'b0;
  assign result_o[32] = 1'b0;
  assign result_o[33] = 1'b0;
  assign result_o[34] = 1'b0;
  assign result_o[35] = 1'b0;
  assign result_o[36] = 1'b0;
  assign result_o[37] = 1'b0;
  assign result_o[38] = 1'b0;
  assign result_o[39] = 1'b0;
  assign result_o[40] = 1'b0;
  assign result_o[41] = 1'b0;
  assign result_o[42] = 1'b0;
  assign result_o[43] = 1'b0;
  assign result_o[44] = 1'b0;
  assign result_o[45] = 1'b0;
  assign result_o[46] = 1'b0;
  assign result_o[47] = 1'b0;
  assign result_o[48] = 1'b0;
  assign result_o[49] = 1'b0;
  assign result_o[50] = 1'b0;
  assign result_o[51] = 1'b0;
  assign result_o[52] = 1'b0;
  assign result_o[53] = 1'b0;
  assign result_o[54] = 1'b0;
  assign result_o[55] = 1'b0;
  assign result_o[56] = 1'b0;
  assign result_o[57] = 1'b0;
  assign result_o[58] = 1'b0;
  assign result_o[59] = 1'b0;
  assign result_o[60] = 1'b0;
  assign result_o[61] = 1'b0;
  assign result_o[62] = 1'b0;
  assign result_o[63] = 1'b0;

endmodule



module bsg_dff_width_p1890
(
  clk_i,
  data_i,
  data_o
);

  input [1889:0] data_i;
  output [1889:0] data_o;
  input clk_i;
  reg [1889:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[1889:0] } <= { data_i[1889:0] };
    end 
  end


endmodule



module bsg_mux_segmented_segments_p5_segment_width_p128
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [639:0] data0_i;
  input [639:0] data1_i;
  input [4:0] sel_i;
  output [639:0] data_o;
  wire [639:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9;
  assign data_o[127:0] = (N0)? data1_i[127:0] : 
                         (N5)? data0_i[127:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[255:128] = (N1)? data1_i[255:128] : 
                           (N6)? data0_i[255:128] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[383:256] = (N2)? data1_i[383:256] : 
                           (N7)? data0_i[383:256] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[511:384] = (N3)? data1_i[511:384] : 
                           (N8)? data0_i[511:384] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[639:512] = (N4)? data1_i[639:512] : 
                           (N9)? data0_i[639:512] : 1'b0;
  assign N4 = sel_i[4];
  assign N5 = ~sel_i[0];
  assign N6 = ~sel_i[1];
  assign N7 = ~sel_i[2];
  assign N8 = ~sel_i[3];
  assign N9 = ~sel_i[4];

endmodule



module bsg_dff_width_p640
(
  clk_i,
  data_i,
  data_o
);

  input [639:0] data_i;
  output [639:0] data_o;
  input clk_i;
  reg [639:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[639:0] } <= { data_i[639:0] };
    end 
  end


endmodule



module bsg_dff_width_p35
(
  clk_i,
  data_i,
  data_o
);

  input [34:0] data_i;
  output [34:0] data_o;
  input clk_i;
  reg [34:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[34:0] } <= { data_i[34:0] };
    end 
  end


endmodule



module bp_be_calculator_top_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_core_els_p1_num_lce_p2_lce_sets_p64_cce_block_size_in_bytes_p64
(
  clk_i,
  reset_i,
  proc_cfg_i,
  issue_pkt_i,
  issue_pkt_v_i,
  issue_pkt_ready_o,
  chk_dispatch_v_i,
  chk_roll_i,
  chk_poison_ex_i,
  chk_poison_isd_i,
  calc_status_o,
  mmu_cmd_o,
  mmu_cmd_v_o,
  mmu_cmd_ready_i,
  mmu_resp_i,
  mmu_resp_v_i,
  mmu_resp_ready_o,
  cmt_trace_stage_reg_o,
  cmt_trace_result_o,
  cmt_trace_exc_o,
  decoded_fu_op_o
);

  input [2:0] proc_cfg_i;
  input [220:0] issue_pkt_i;
  output [301:0] calc_status_o;
  output [123:0] mmu_cmd_o;
  input [70:0] mmu_resp_i;
  output [377:0] cmt_trace_stage_reg_o;
  output [127:0] cmt_trace_result_o;
  output [6:0] cmt_trace_exc_o;
  output [3:0] decoded_fu_op_o;
  input clk_i;
  input reset_i;
  input issue_pkt_v_i;
  input chk_dispatch_v_i;
  input chk_roll_i;
  input chk_poison_ex_i;
  input chk_poison_isd_i;
  input mmu_cmd_ready_i;
  input mmu_resp_v_i;
  output issue_pkt_ready_o;
  output mmu_cmd_v_o;
  output mmu_resp_ready_o;
  wire [301:0] calc_status_o;
  wire [123:0] mmu_cmd_o;
  wire [377:0] cmt_trace_stage_reg_o;
  wire [127:0] cmt_trace_result_o,mul_calc_result,mem_calc_result,fp_calc_result,
  nop_calc_result;
  wire [6:0] cmt_trace_exc_o;
  wire [3:0] decoded_fu_op_o;
  wire issue_pkt_ready_o,mmu_cmd_v_o,mmu_resp_ready_o,decoded_fp_not_int_v_,
  decoded_rs1_addr__4_,decoded_rs1_addr__3_,decoded_rs1_addr__2_,decoded_rs1_addr__1_,
  decoded_rs1_addr__0_,decoded_rs2_addr__4_,decoded_rs2_addr__3_,decoded_rs2_addr__2_,
  decoded_rs2_addr__1_,decoded_rs2_addr__0_,n_0_net_,comp_stage_r_3__result__63_,
  comp_stage_r_3__result__62_,comp_stage_r_3__result__61_,comp_stage_r_3__result__60_,
  comp_stage_r_3__result__59_,comp_stage_r_3__result__58_,
  comp_stage_r_3__result__57_,comp_stage_r_3__result__56_,comp_stage_r_3__result__55_,
  comp_stage_r_3__result__54_,comp_stage_r_3__result__53_,comp_stage_r_3__result__52_,
  comp_stage_r_3__result__51_,comp_stage_r_3__result__50_,comp_stage_r_3__result__49_,
  comp_stage_r_3__result__48_,comp_stage_r_3__result__47_,comp_stage_r_3__result__46_,
  comp_stage_r_3__result__45_,comp_stage_r_3__result__44_,comp_stage_r_3__result__43_,
  comp_stage_r_3__result__42_,comp_stage_r_3__result__41_,comp_stage_r_3__result__40_,
  comp_stage_r_3__result__39_,comp_stage_r_3__result__38_,
  comp_stage_r_3__result__37_,comp_stage_r_3__result__36_,comp_stage_r_3__result__35_,
  comp_stage_r_3__result__34_,comp_stage_r_3__result__33_,comp_stage_r_3__result__32_,
  comp_stage_r_3__result__31_,comp_stage_r_3__result__30_,comp_stage_r_3__result__29_,
  comp_stage_r_3__result__28_,comp_stage_r_3__result__27_,comp_stage_r_3__result__26_,
  comp_stage_r_3__result__25_,comp_stage_r_3__result__24_,comp_stage_r_3__result__23_,
  comp_stage_r_3__result__22_,comp_stage_r_3__result__21_,comp_stage_r_3__result__20_,
  comp_stage_r_3__result__19_,comp_stage_r_3__result__18_,
  comp_stage_r_3__result__17_,comp_stage_r_3__result__16_,comp_stage_r_3__result__15_,
  comp_stage_r_3__result__14_,comp_stage_r_3__result__13_,comp_stage_r_3__result__12_,
  comp_stage_r_3__result__11_,comp_stage_r_3__result__10_,comp_stage_r_3__result__9_,
  comp_stage_r_3__result__8_,comp_stage_r_3__result__7_,comp_stage_r_3__result__6_,
  comp_stage_r_3__result__5_,comp_stage_r_3__result__4_,comp_stage_r_3__result__3_,
  comp_stage_r_3__result__2_,comp_stage_r_3__result__1_,comp_stage_r_3__result__0_,
  comp_stage_r_3__br_tgt__63_,comp_stage_r_3__br_tgt__62_,comp_stage_r_3__br_tgt__61_,
  comp_stage_r_3__br_tgt__60_,comp_stage_r_3__br_tgt__59_,comp_stage_r_3__br_tgt__58_,
  comp_stage_r_3__br_tgt__57_,comp_stage_r_3__br_tgt__56_,
  comp_stage_r_3__br_tgt__55_,comp_stage_r_3__br_tgt__54_,comp_stage_r_3__br_tgt__53_,
  comp_stage_r_3__br_tgt__52_,comp_stage_r_3__br_tgt__51_,comp_stage_r_3__br_tgt__50_,
  comp_stage_r_3__br_tgt__49_,comp_stage_r_3__br_tgt__48_,comp_stage_r_3__br_tgt__47_,
  comp_stage_r_3__br_tgt__46_,comp_stage_r_3__br_tgt__45_,comp_stage_r_3__br_tgt__44_,
  comp_stage_r_3__br_tgt__43_,comp_stage_r_3__br_tgt__42_,comp_stage_r_3__br_tgt__41_,
  comp_stage_r_3__br_tgt__40_,comp_stage_r_3__br_tgt__39_,comp_stage_r_3__br_tgt__38_,
  comp_stage_r_3__br_tgt__37_,comp_stage_r_3__br_tgt__36_,
  comp_stage_r_3__br_tgt__35_,comp_stage_r_3__br_tgt__34_,comp_stage_r_3__br_tgt__33_,
  comp_stage_r_3__br_tgt__32_,comp_stage_r_3__br_tgt__31_,comp_stage_r_3__br_tgt__30_,
  comp_stage_r_3__br_tgt__29_,comp_stage_r_3__br_tgt__28_,comp_stage_r_3__br_tgt__27_,
  comp_stage_r_3__br_tgt__26_,comp_stage_r_3__br_tgt__25_,comp_stage_r_3__br_tgt__24_,
  comp_stage_r_3__br_tgt__23_,comp_stage_r_3__br_tgt__22_,comp_stage_r_3__br_tgt__21_,
  comp_stage_r_3__br_tgt__20_,comp_stage_r_3__br_tgt__19_,comp_stage_r_3__br_tgt__18_,
  comp_stage_r_3__br_tgt__17_,comp_stage_r_3__br_tgt__16_,
  comp_stage_r_3__br_tgt__15_,comp_stage_r_3__br_tgt__14_,comp_stage_r_3__br_tgt__13_,
  comp_stage_r_3__br_tgt__12_,comp_stage_r_3__br_tgt__11_,comp_stage_r_3__br_tgt__10_,
  comp_stage_r_3__br_tgt__9_,comp_stage_r_3__br_tgt__8_,comp_stage_r_3__br_tgt__7_,
  comp_stage_r_3__br_tgt__6_,comp_stage_r_3__br_tgt__5_,comp_stage_r_3__br_tgt__4_,
  comp_stage_r_3__br_tgt__3_,comp_stage_r_3__br_tgt__2_,comp_stage_r_3__br_tgt__1_,
  comp_stage_r_3__br_tgt__0_,comp_stage_r_2__result__63_,comp_stage_r_2__result__62_,
  comp_stage_r_2__result__61_,comp_stage_r_2__result__60_,comp_stage_r_2__result__59_,
  comp_stage_r_2__result__58_,comp_stage_r_2__result__57_,comp_stage_r_2__result__56_,
  comp_stage_r_2__result__55_,comp_stage_r_2__result__54_,comp_stage_r_2__result__53_,
  comp_stage_r_2__result__52_,comp_stage_r_2__result__51_,
  comp_stage_r_2__result__50_,comp_stage_r_2__result__49_,comp_stage_r_2__result__48_,
  comp_stage_r_2__result__47_,comp_stage_r_2__result__46_,comp_stage_r_2__result__45_,
  comp_stage_r_2__result__44_,comp_stage_r_2__result__43_,comp_stage_r_2__result__42_,
  comp_stage_r_2__result__41_,comp_stage_r_2__result__40_,comp_stage_r_2__result__39_,
  comp_stage_r_2__result__38_,comp_stage_r_2__result__37_,comp_stage_r_2__result__36_,
  comp_stage_r_2__result__35_,comp_stage_r_2__result__34_,comp_stage_r_2__result__33_,
  comp_stage_r_2__result__32_,comp_stage_r_2__result__31_,
  comp_stage_r_2__result__30_,comp_stage_r_2__result__29_,comp_stage_r_2__result__28_,
  comp_stage_r_2__result__27_,comp_stage_r_2__result__26_,comp_stage_r_2__result__25_,
  comp_stage_r_2__result__24_,comp_stage_r_2__result__23_,comp_stage_r_2__result__22_,
  comp_stage_r_2__result__21_,comp_stage_r_2__result__20_,comp_stage_r_2__result__19_,
  comp_stage_r_2__result__18_,comp_stage_r_2__result__17_,comp_stage_r_2__result__16_,
  comp_stage_r_2__result__15_,comp_stage_r_2__result__14_,comp_stage_r_2__result__13_,
  comp_stage_r_2__result__12_,comp_stage_r_2__result__11_,
  comp_stage_r_2__result__10_,comp_stage_r_2__result__9_,comp_stage_r_2__result__8_,
  comp_stage_r_2__result__7_,comp_stage_r_2__result__6_,comp_stage_r_2__result__5_,
  comp_stage_r_2__result__4_,comp_stage_r_2__result__3_,comp_stage_r_2__result__2_,
  comp_stage_r_2__result__1_,comp_stage_r_2__result__0_,comp_stage_r_2__br_tgt__63_,
  comp_stage_r_2__br_tgt__62_,comp_stage_r_2__br_tgt__61_,comp_stage_r_2__br_tgt__60_,
  comp_stage_r_2__br_tgt__59_,comp_stage_r_2__br_tgt__58_,comp_stage_r_2__br_tgt__57_,
  comp_stage_r_2__br_tgt__56_,comp_stage_r_2__br_tgt__55_,comp_stage_r_2__br_tgt__54_,
  comp_stage_r_2__br_tgt__53_,comp_stage_r_2__br_tgt__52_,comp_stage_r_2__br_tgt__51_,
  comp_stage_r_2__br_tgt__50_,comp_stage_r_2__br_tgt__49_,
  comp_stage_r_2__br_tgt__48_,comp_stage_r_2__br_tgt__47_,comp_stage_r_2__br_tgt__46_,
  comp_stage_r_2__br_tgt__45_,comp_stage_r_2__br_tgt__44_,comp_stage_r_2__br_tgt__43_,
  comp_stage_r_2__br_tgt__42_,comp_stage_r_2__br_tgt__41_,comp_stage_r_2__br_tgt__40_,
  comp_stage_r_2__br_tgt__39_,comp_stage_r_2__br_tgt__38_,comp_stage_r_2__br_tgt__37_,
  comp_stage_r_2__br_tgt__36_,comp_stage_r_2__br_tgt__35_,comp_stage_r_2__br_tgt__34_,
  comp_stage_r_2__br_tgt__33_,comp_stage_r_2__br_tgt__32_,comp_stage_r_2__br_tgt__31_,
  comp_stage_r_2__br_tgt__30_,comp_stage_r_2__br_tgt__29_,
  comp_stage_r_2__br_tgt__28_,comp_stage_r_2__br_tgt__27_,comp_stage_r_2__br_tgt__26_,
  comp_stage_r_2__br_tgt__25_,comp_stage_r_2__br_tgt__24_,comp_stage_r_2__br_tgt__23_,
  comp_stage_r_2__br_tgt__22_,comp_stage_r_2__br_tgt__21_,comp_stage_r_2__br_tgt__20_,
  comp_stage_r_2__br_tgt__19_,comp_stage_r_2__br_tgt__18_,comp_stage_r_2__br_tgt__17_,
  comp_stage_r_2__br_tgt__16_,comp_stage_r_2__br_tgt__15_,comp_stage_r_2__br_tgt__14_,
  comp_stage_r_2__br_tgt__13_,comp_stage_r_2__br_tgt__12_,comp_stage_r_2__br_tgt__11_,
  comp_stage_r_2__br_tgt__10_,comp_stage_r_2__br_tgt__9_,comp_stage_r_2__br_tgt__8_,
  comp_stage_r_2__br_tgt__7_,comp_stage_r_2__br_tgt__6_,
  comp_stage_r_2__br_tgt__5_,comp_stage_r_2__br_tgt__4_,comp_stage_r_2__br_tgt__3_,
  comp_stage_r_2__br_tgt__2_,comp_stage_r_2__br_tgt__1_,comp_stage_r_2__br_tgt__0_,
  comp_stage_r_1__result__63_,comp_stage_r_1__result__62_,comp_stage_r_1__result__61_,
  comp_stage_r_1__result__60_,comp_stage_r_1__result__59_,comp_stage_r_1__result__58_,
  comp_stage_r_1__result__57_,comp_stage_r_1__result__56_,comp_stage_r_1__result__55_,
  comp_stage_r_1__result__54_,comp_stage_r_1__result__53_,comp_stage_r_1__result__52_,
  comp_stage_r_1__result__51_,comp_stage_r_1__result__50_,comp_stage_r_1__result__49_,
  comp_stage_r_1__result__48_,comp_stage_r_1__result__47_,comp_stage_r_1__result__46_,
  comp_stage_r_1__result__45_,comp_stage_r_1__result__44_,
  comp_stage_r_1__result__43_,comp_stage_r_1__result__42_,comp_stage_r_1__result__41_,
  comp_stage_r_1__result__40_,comp_stage_r_1__result__39_,comp_stage_r_1__result__38_,
  comp_stage_r_1__result__37_,comp_stage_r_1__result__36_,comp_stage_r_1__result__35_,
  comp_stage_r_1__result__34_,comp_stage_r_1__result__33_,comp_stage_r_1__result__32_,
  comp_stage_r_1__result__31_,comp_stage_r_1__result__30_,comp_stage_r_1__result__29_,
  comp_stage_r_1__result__28_,comp_stage_r_1__result__27_,comp_stage_r_1__result__26_,
  comp_stage_r_1__result__25_,comp_stage_r_1__result__24_,
  comp_stage_r_1__result__23_,comp_stage_r_1__result__22_,comp_stage_r_1__result__21_,
  comp_stage_r_1__result__20_,comp_stage_r_1__result__19_,comp_stage_r_1__result__18_,
  comp_stage_r_1__result__17_,comp_stage_r_1__result__16_,comp_stage_r_1__result__15_,
  comp_stage_r_1__result__14_,comp_stage_r_1__result__13_,comp_stage_r_1__result__12_,
  comp_stage_r_1__result__11_,comp_stage_r_1__result__10_,comp_stage_r_1__result__9_,
  comp_stage_r_1__result__8_,comp_stage_r_1__result__7_,comp_stage_r_1__result__6_,
  comp_stage_r_1__result__5_,comp_stage_r_1__result__4_,comp_stage_r_1__result__3_,
  comp_stage_r_1__result__2_,comp_stage_r_1__result__1_,comp_stage_r_1__result__0_,
  comp_stage_r_1__br_tgt__63_,comp_stage_r_1__br_tgt__62_,
  comp_stage_r_1__br_tgt__61_,comp_stage_r_1__br_tgt__60_,comp_stage_r_1__br_tgt__59_,
  comp_stage_r_1__br_tgt__58_,comp_stage_r_1__br_tgt__57_,comp_stage_r_1__br_tgt__56_,
  comp_stage_r_1__br_tgt__55_,comp_stage_r_1__br_tgt__54_,comp_stage_r_1__br_tgt__53_,
  comp_stage_r_1__br_tgt__52_,comp_stage_r_1__br_tgt__51_,comp_stage_r_1__br_tgt__50_,
  comp_stage_r_1__br_tgt__49_,comp_stage_r_1__br_tgt__48_,comp_stage_r_1__br_tgt__47_,
  comp_stage_r_1__br_tgt__46_,comp_stage_r_1__br_tgt__45_,comp_stage_r_1__br_tgt__44_,
  comp_stage_r_1__br_tgt__43_,comp_stage_r_1__br_tgt__42_,
  comp_stage_r_1__br_tgt__41_,comp_stage_r_1__br_tgt__40_,comp_stage_r_1__br_tgt__39_,
  comp_stage_r_1__br_tgt__38_,comp_stage_r_1__br_tgt__37_,comp_stage_r_1__br_tgt__36_,
  comp_stage_r_1__br_tgt__35_,comp_stage_r_1__br_tgt__34_,comp_stage_r_1__br_tgt__33_,
  comp_stage_r_1__br_tgt__32_,comp_stage_r_1__br_tgt__31_,comp_stage_r_1__br_tgt__30_,
  comp_stage_r_1__br_tgt__29_,comp_stage_r_1__br_tgt__28_,comp_stage_r_1__br_tgt__27_,
  comp_stage_r_1__br_tgt__26_,comp_stage_r_1__br_tgt__25_,comp_stage_r_1__br_tgt__24_,
  comp_stage_r_1__br_tgt__23_,comp_stage_r_1__br_tgt__22_,
  comp_stage_r_1__br_tgt__21_,comp_stage_r_1__br_tgt__20_,comp_stage_r_1__br_tgt__19_,
  comp_stage_r_1__br_tgt__18_,comp_stage_r_1__br_tgt__17_,comp_stage_r_1__br_tgt__16_,
  comp_stage_r_1__br_tgt__15_,comp_stage_r_1__br_tgt__14_,comp_stage_r_1__br_tgt__13_,
  comp_stage_r_1__br_tgt__12_,comp_stage_r_1__br_tgt__11_,comp_stage_r_1__br_tgt__10_,
  comp_stage_r_1__br_tgt__9_,comp_stage_r_1__br_tgt__8_,comp_stage_r_1__br_tgt__7_,
  comp_stage_r_1__br_tgt__6_,comp_stage_r_1__br_tgt__5_,comp_stage_r_1__br_tgt__4_,
  comp_stage_r_1__br_tgt__3_,comp_stage_r_1__br_tgt__2_,comp_stage_r_1__br_tgt__1_,
  comp_stage_r_1__br_tgt__0_,comp_stage_r_0__result__63_,comp_stage_r_0__result__62_,
  comp_stage_r_0__result__61_,comp_stage_r_0__result__60_,comp_stage_r_0__result__59_,
  comp_stage_r_0__result__58_,comp_stage_r_0__result__57_,
  comp_stage_r_0__result__56_,comp_stage_r_0__result__55_,comp_stage_r_0__result__54_,
  comp_stage_r_0__result__53_,comp_stage_r_0__result__52_,comp_stage_r_0__result__51_,
  comp_stage_r_0__result__50_,comp_stage_r_0__result__49_,comp_stage_r_0__result__48_,
  comp_stage_r_0__result__47_,comp_stage_r_0__result__46_,comp_stage_r_0__result__45_,
  comp_stage_r_0__result__44_,comp_stage_r_0__result__43_,comp_stage_r_0__result__42_,
  comp_stage_r_0__result__41_,comp_stage_r_0__result__40_,comp_stage_r_0__result__39_,
  comp_stage_r_0__result__38_,comp_stage_r_0__result__37_,
  comp_stage_r_0__result__36_,comp_stage_r_0__result__35_,comp_stage_r_0__result__34_,
  comp_stage_r_0__result__33_,comp_stage_r_0__result__32_,comp_stage_r_0__result__31_,
  comp_stage_r_0__result__30_,comp_stage_r_0__result__29_,comp_stage_r_0__result__28_,
  comp_stage_r_0__result__27_,comp_stage_r_0__result__26_,comp_stage_r_0__result__25_,
  comp_stage_r_0__result__24_,comp_stage_r_0__result__23_,comp_stage_r_0__result__22_,
  comp_stage_r_0__result__21_,comp_stage_r_0__result__20_,comp_stage_r_0__result__19_,
  comp_stage_r_0__result__18_,comp_stage_r_0__result__17_,
  comp_stage_r_0__result__16_,comp_stage_r_0__result__15_,comp_stage_r_0__result__14_,
  comp_stage_r_0__result__13_,comp_stage_r_0__result__12_,comp_stage_r_0__result__11_,
  comp_stage_r_0__result__10_,comp_stage_r_0__result__9_,comp_stage_r_0__result__8_,
  comp_stage_r_0__result__7_,comp_stage_r_0__result__6_,comp_stage_r_0__result__5_,
  comp_stage_r_0__result__4_,comp_stage_r_0__result__3_,comp_stage_r_0__result__2_,
  comp_stage_r_0__result__1_,comp_stage_r_0__result__0_,comp_stage_r_0__br_tgt__63_,
  comp_stage_r_0__br_tgt__62_,comp_stage_r_0__br_tgt__61_,comp_stage_r_0__br_tgt__60_,
  comp_stage_r_0__br_tgt__59_,comp_stage_r_0__br_tgt__58_,comp_stage_r_0__br_tgt__57_,
  comp_stage_r_0__br_tgt__56_,comp_stage_r_0__br_tgt__55_,
  comp_stage_r_0__br_tgt__54_,comp_stage_r_0__br_tgt__53_,comp_stage_r_0__br_tgt__52_,
  comp_stage_r_0__br_tgt__51_,comp_stage_r_0__br_tgt__50_,comp_stage_r_0__br_tgt__49_,
  comp_stage_r_0__br_tgt__48_,comp_stage_r_0__br_tgt__47_,comp_stage_r_0__br_tgt__46_,
  comp_stage_r_0__br_tgt__45_,comp_stage_r_0__br_tgt__44_,comp_stage_r_0__br_tgt__43_,
  comp_stage_r_0__br_tgt__42_,comp_stage_r_0__br_tgt__41_,comp_stage_r_0__br_tgt__40_,
  comp_stage_r_0__br_tgt__39_,comp_stage_r_0__br_tgt__38_,comp_stage_r_0__br_tgt__37_,
  comp_stage_r_0__br_tgt__36_,comp_stage_r_0__br_tgt__35_,
  comp_stage_r_0__br_tgt__34_,comp_stage_r_0__br_tgt__33_,comp_stage_r_0__br_tgt__32_,
  comp_stage_r_0__br_tgt__31_,comp_stage_r_0__br_tgt__30_,comp_stage_r_0__br_tgt__29_,
  comp_stage_r_0__br_tgt__28_,comp_stage_r_0__br_tgt__27_,comp_stage_r_0__br_tgt__26_,
  comp_stage_r_0__br_tgt__25_,comp_stage_r_0__br_tgt__24_,comp_stage_r_0__br_tgt__23_,
  comp_stage_r_0__br_tgt__22_,comp_stage_r_0__br_tgt__21_,comp_stage_r_0__br_tgt__20_,
  comp_stage_r_0__br_tgt__19_,comp_stage_r_0__br_tgt__18_,comp_stage_r_0__br_tgt__17_,
  comp_stage_r_0__br_tgt__16_,comp_stage_r_0__br_tgt__15_,
  comp_stage_r_0__br_tgt__14_,comp_stage_r_0__br_tgt__13_,comp_stage_r_0__br_tgt__12_,
  comp_stage_r_0__br_tgt__11_,comp_stage_r_0__br_tgt__10_,comp_stage_r_0__br_tgt__9_,
  comp_stage_r_0__br_tgt__8_,comp_stage_r_0__br_tgt__7_,comp_stage_r_0__br_tgt__6_,
  comp_stage_r_0__br_tgt__5_,comp_stage_r_0__br_tgt__4_,comp_stage_r_0__br_tgt__3_,
  comp_stage_r_0__br_tgt__2_,comp_stage_r_0__br_tgt__1_,comp_stage_r_0__br_tgt__0_,
  calc_stage_r_3__instr_metadata__itag__7_,calc_stage_r_3__instr_metadata__itag__6_,
  calc_stage_r_3__instr_metadata__itag__5_,calc_stage_r_3__instr_metadata__itag__4_,
  calc_stage_r_3__instr_metadata__itag__3_,calc_stage_r_3__instr_metadata__itag__2_,
  calc_stage_r_3__instr_metadata__itag__1_,calc_stage_r_3__instr_metadata__itag__0_,
  calc_stage_r_3__instr_metadata__pc__63_,calc_stage_r_3__instr_metadata__pc__62_,
  calc_stage_r_3__instr_metadata__pc__61_,calc_stage_r_3__instr_metadata__pc__60_,
  calc_stage_r_3__instr_metadata__pc__59_,calc_stage_r_3__instr_metadata__pc__58_,
  calc_stage_r_3__instr_metadata__pc__57_,calc_stage_r_3__instr_metadata__pc__56_,
  calc_stage_r_3__instr_metadata__pc__55_,calc_stage_r_3__instr_metadata__pc__54_,
  calc_stage_r_3__instr_metadata__pc__53_,calc_stage_r_3__instr_metadata__pc__52_,
  calc_stage_r_3__instr_metadata__pc__51_,calc_stage_r_3__instr_metadata__pc__50_,
  calc_stage_r_3__instr_metadata__pc__49_,calc_stage_r_3__instr_metadata__pc__48_,
  calc_stage_r_3__instr_metadata__pc__47_,calc_stage_r_3__instr_metadata__pc__46_,
  calc_stage_r_3__instr_metadata__pc__45_,calc_stage_r_3__instr_metadata__pc__44_,
  calc_stage_r_3__instr_metadata__pc__43_,calc_stage_r_3__instr_metadata__pc__42_,
  calc_stage_r_3__instr_metadata__pc__41_,calc_stage_r_3__instr_metadata__pc__40_,
  calc_stage_r_3__instr_metadata__pc__39_,calc_stage_r_3__instr_metadata__pc__38_,
  calc_stage_r_3__instr_metadata__pc__37_,calc_stage_r_3__instr_metadata__pc__36_,
  calc_stage_r_3__instr_metadata__pc__35_,calc_stage_r_3__instr_metadata__pc__34_,
  calc_stage_r_3__instr_metadata__pc__33_,calc_stage_r_3__instr_metadata__pc__32_,
  calc_stage_r_3__instr_metadata__pc__31_,calc_stage_r_3__instr_metadata__pc__30_,
  calc_stage_r_3__instr_metadata__pc__29_,calc_stage_r_3__instr_metadata__pc__28_,
  calc_stage_r_3__instr_metadata__pc__27_,calc_stage_r_3__instr_metadata__pc__26_,
  calc_stage_r_3__instr_metadata__pc__25_,calc_stage_r_3__instr_metadata__pc__24_,
  calc_stage_r_3__instr_metadata__pc__23_,calc_stage_r_3__instr_metadata__pc__22_,
  calc_stage_r_3__instr_metadata__pc__21_,calc_stage_r_3__instr_metadata__pc__20_,
  calc_stage_r_3__instr_metadata__pc__19_,calc_stage_r_3__instr_metadata__pc__18_,
  calc_stage_r_3__instr_metadata__pc__17_,calc_stage_r_3__instr_metadata__pc__16_,
  calc_stage_r_3__instr_metadata__pc__15_,calc_stage_r_3__instr_metadata__pc__14_,
  calc_stage_r_3__instr_metadata__pc__13_,calc_stage_r_3__instr_metadata__pc__12_,
  calc_stage_r_3__instr_metadata__pc__11_,calc_stage_r_3__instr_metadata__pc__10_,
  calc_stage_r_3__instr_metadata__pc__9_,calc_stage_r_3__instr_metadata__pc__8_,
  calc_stage_r_3__instr_metadata__pc__7_,calc_stage_r_3__instr_metadata__pc__6_,
  calc_stage_r_3__instr_metadata__pc__5_,calc_stage_r_3__instr_metadata__pc__4_,
  calc_stage_r_3__instr_metadata__pc__3_,calc_stage_r_3__instr_metadata__pc__2_,
  calc_stage_r_3__instr_metadata__pc__1_,calc_stage_r_3__instr_metadata__pc__0_,
  calc_stage_r_3__instr_metadata__fe_exception_not_instr_,
  calc_stage_r_3__instr_metadata__fe_exception_code__1_,calc_stage_r_3__instr_metadata__fe_exception_code__0_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__35_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__34_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__33_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__32_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__31_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__30_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__29_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__28_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__27_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__26_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__25_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__24_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__23_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__22_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__21_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__20_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__19_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__18_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__17_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__16_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__15_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__14_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__13_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__12_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__11_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__10_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__9_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__8_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__7_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__6_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__5_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__4_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__3_,calc_stage_r_3__instr_metadata__branch_metadata_fwd__2_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__1_,
  calc_stage_r_3__instr_metadata__branch_metadata_fwd__0_,calc_stage_r_3__instr__31_,
  calc_stage_r_3__instr__30_,calc_stage_r_3__instr__29_,calc_stage_r_3__instr__28_,
  calc_stage_r_3__instr__27_,calc_stage_r_3__instr__26_,calc_stage_r_3__instr__25_,
  calc_stage_r_3__instr__24_,calc_stage_r_3__instr__23_,calc_stage_r_3__instr__22_,
  calc_stage_r_3__instr__21_,calc_stage_r_3__instr__20_,calc_stage_r_3__instr__19_,
  calc_stage_r_3__instr__18_,calc_stage_r_3__instr__17_,calc_stage_r_3__instr__16_,
  calc_stage_r_3__instr__15_,calc_stage_r_3__instr__14_,calc_stage_r_3__instr__13_,
  calc_stage_r_3__instr__12_,calc_stage_r_3__instr__11_,calc_stage_r_3__instr__10_,
  calc_stage_r_3__instr__9_,calc_stage_r_3__instr__8_,calc_stage_r_3__instr__7_,
  calc_stage_r_3__instr__6_,calc_stage_r_3__instr__5_,calc_stage_r_3__instr__4_,
  calc_stage_r_3__instr__3_,calc_stage_r_3__instr__2_,calc_stage_r_3__instr__1_,
  calc_stage_r_3__instr__0_,calc_stage_r_3__instr_operands__rs1__63_,
  calc_stage_r_3__instr_operands__rs1__62_,calc_stage_r_3__instr_operands__rs1__61_,
  calc_stage_r_3__instr_operands__rs1__60_,calc_stage_r_3__instr_operands__rs1__59_,
  calc_stage_r_3__instr_operands__rs1__58_,calc_stage_r_3__instr_operands__rs1__57_,
  calc_stage_r_3__instr_operands__rs1__56_,calc_stage_r_3__instr_operands__rs1__55_,
  calc_stage_r_3__instr_operands__rs1__54_,calc_stage_r_3__instr_operands__rs1__53_,
  calc_stage_r_3__instr_operands__rs1__52_,calc_stage_r_3__instr_operands__rs1__51_,
  calc_stage_r_3__instr_operands__rs1__50_,calc_stage_r_3__instr_operands__rs1__49_,
  calc_stage_r_3__instr_operands__rs1__48_,calc_stage_r_3__instr_operands__rs1__47_,
  calc_stage_r_3__instr_operands__rs1__46_,calc_stage_r_3__instr_operands__rs1__45_,
  calc_stage_r_3__instr_operands__rs1__44_,calc_stage_r_3__instr_operands__rs1__43_,
  calc_stage_r_3__instr_operands__rs1__42_,calc_stage_r_3__instr_operands__rs1__41_,
  calc_stage_r_3__instr_operands__rs1__40_,calc_stage_r_3__instr_operands__rs1__39_,
  calc_stage_r_3__instr_operands__rs1__38_,calc_stage_r_3__instr_operands__rs1__37_,
  calc_stage_r_3__instr_operands__rs1__36_,calc_stage_r_3__instr_operands__rs1__35_,
  calc_stage_r_3__instr_operands__rs1__34_,calc_stage_r_3__instr_operands__rs1__33_,
  calc_stage_r_3__instr_operands__rs1__32_,calc_stage_r_3__instr_operands__rs1__31_,
  calc_stage_r_3__instr_operands__rs1__30_,calc_stage_r_3__instr_operands__rs1__29_,
  calc_stage_r_3__instr_operands__rs1__28_,calc_stage_r_3__instr_operands__rs1__27_,
  calc_stage_r_3__instr_operands__rs1__26_,
  calc_stage_r_3__instr_operands__rs1__25_,calc_stage_r_3__instr_operands__rs1__24_,
  calc_stage_r_3__instr_operands__rs1__23_,calc_stage_r_3__instr_operands__rs1__22_,
  calc_stage_r_3__instr_operands__rs1__21_,calc_stage_r_3__instr_operands__rs1__20_,
  calc_stage_r_3__instr_operands__rs1__19_,calc_stage_r_3__instr_operands__rs1__18_,
  calc_stage_r_3__instr_operands__rs1__17_,calc_stage_r_3__instr_operands__rs1__16_,
  calc_stage_r_3__instr_operands__rs1__15_,calc_stage_r_3__instr_operands__rs1__14_,
  calc_stage_r_3__instr_operands__rs1__13_,calc_stage_r_3__instr_operands__rs1__12_,
  calc_stage_r_3__instr_operands__rs1__11_,calc_stage_r_3__instr_operands__rs1__10_,
  calc_stage_r_3__instr_operands__rs1__9_,calc_stage_r_3__instr_operands__rs1__8_,
  calc_stage_r_3__instr_operands__rs1__7_,calc_stage_r_3__instr_operands__rs1__6_,
  calc_stage_r_3__instr_operands__rs1__5_,calc_stage_r_3__instr_operands__rs1__4_,
  calc_stage_r_3__instr_operands__rs1__3_,calc_stage_r_3__instr_operands__rs1__2_,
  calc_stage_r_3__instr_operands__rs1__1_,calc_stage_r_3__instr_operands__rs1__0_,
  calc_stage_r_3__instr_operands__rs2__63_,calc_stage_r_3__instr_operands__rs2__62_,
  calc_stage_r_3__instr_operands__rs2__61_,calc_stage_r_3__instr_operands__rs2__60_,
  calc_stage_r_3__instr_operands__rs2__59_,calc_stage_r_3__instr_operands__rs2__58_,
  calc_stage_r_3__instr_operands__rs2__57_,calc_stage_r_3__instr_operands__rs2__56_,
  calc_stage_r_3__instr_operands__rs2__55_,calc_stage_r_3__instr_operands__rs2__54_,
  calc_stage_r_3__instr_operands__rs2__53_,calc_stage_r_3__instr_operands__rs2__52_,
  calc_stage_r_3__instr_operands__rs2__51_,calc_stage_r_3__instr_operands__rs2__50_,
  calc_stage_r_3__instr_operands__rs2__49_,calc_stage_r_3__instr_operands__rs2__48_,
  calc_stage_r_3__instr_operands__rs2__47_,calc_stage_r_3__instr_operands__rs2__46_,
  calc_stage_r_3__instr_operands__rs2__45_,calc_stage_r_3__instr_operands__rs2__44_,
  calc_stage_r_3__instr_operands__rs2__43_,calc_stage_r_3__instr_operands__rs2__42_,
  calc_stage_r_3__instr_operands__rs2__41_,calc_stage_r_3__instr_operands__rs2__40_,
  calc_stage_r_3__instr_operands__rs2__39_,
  calc_stage_r_3__instr_operands__rs2__38_,calc_stage_r_3__instr_operands__rs2__37_,
  calc_stage_r_3__instr_operands__rs2__36_,calc_stage_r_3__instr_operands__rs2__35_,
  calc_stage_r_3__instr_operands__rs2__34_,calc_stage_r_3__instr_operands__rs2__33_,
  calc_stage_r_3__instr_operands__rs2__32_,calc_stage_r_3__instr_operands__rs2__31_,
  calc_stage_r_3__instr_operands__rs2__30_,calc_stage_r_3__instr_operands__rs2__29_,
  calc_stage_r_3__instr_operands__rs2__28_,calc_stage_r_3__instr_operands__rs2__27_,
  calc_stage_r_3__instr_operands__rs2__26_,calc_stage_r_3__instr_operands__rs2__25_,
  calc_stage_r_3__instr_operands__rs2__24_,calc_stage_r_3__instr_operands__rs2__23_,
  calc_stage_r_3__instr_operands__rs2__22_,calc_stage_r_3__instr_operands__rs2__21_,
  calc_stage_r_3__instr_operands__rs2__20_,calc_stage_r_3__instr_operands__rs2__19_,
  calc_stage_r_3__instr_operands__rs2__18_,calc_stage_r_3__instr_operands__rs2__17_,
  calc_stage_r_3__instr_operands__rs2__16_,calc_stage_r_3__instr_operands__rs2__15_,
  calc_stage_r_3__instr_operands__rs2__14_,calc_stage_r_3__instr_operands__rs2__13_,
  calc_stage_r_3__instr_operands__rs2__12_,calc_stage_r_3__instr_operands__rs2__11_,
  calc_stage_r_3__instr_operands__rs2__10_,calc_stage_r_3__instr_operands__rs2__9_,
  calc_stage_r_3__instr_operands__rs2__8_,calc_stage_r_3__instr_operands__rs2__7_,
  calc_stage_r_3__instr_operands__rs2__6_,calc_stage_r_3__instr_operands__rs2__5_,
  calc_stage_r_3__instr_operands__rs2__4_,calc_stage_r_3__instr_operands__rs2__3_,
  calc_stage_r_3__instr_operands__rs2__2_,calc_stage_r_3__instr_operands__rs2__1_,
  calc_stage_r_3__instr_operands__rs2__0_,calc_stage_r_3__instr_operands__imm__63_,
  calc_stage_r_3__instr_operands__imm__62_,calc_stage_r_3__instr_operands__imm__61_,
  calc_stage_r_3__instr_operands__imm__60_,calc_stage_r_3__instr_operands__imm__59_,
  calc_stage_r_3__instr_operands__imm__58_,calc_stage_r_3__instr_operands__imm__57_,
  calc_stage_r_3__instr_operands__imm__56_,calc_stage_r_3__instr_operands__imm__55_,
  calc_stage_r_3__instr_operands__imm__54_,
  calc_stage_r_3__instr_operands__imm__53_,calc_stage_r_3__instr_operands__imm__52_,
  calc_stage_r_3__instr_operands__imm__51_,calc_stage_r_3__instr_operands__imm__50_,
  calc_stage_r_3__instr_operands__imm__49_,calc_stage_r_3__instr_operands__imm__48_,
  calc_stage_r_3__instr_operands__imm__47_,calc_stage_r_3__instr_operands__imm__46_,
  calc_stage_r_3__instr_operands__imm__45_,calc_stage_r_3__instr_operands__imm__44_,
  calc_stage_r_3__instr_operands__imm__43_,calc_stage_r_3__instr_operands__imm__42_,
  calc_stage_r_3__instr_operands__imm__41_,calc_stage_r_3__instr_operands__imm__40_,
  calc_stage_r_3__instr_operands__imm__39_,calc_stage_r_3__instr_operands__imm__38_,
  calc_stage_r_3__instr_operands__imm__37_,calc_stage_r_3__instr_operands__imm__36_,
  calc_stage_r_3__instr_operands__imm__35_,calc_stage_r_3__instr_operands__imm__34_,
  calc_stage_r_3__instr_operands__imm__33_,calc_stage_r_3__instr_operands__imm__32_,
  calc_stage_r_3__instr_operands__imm__31_,calc_stage_r_3__instr_operands__imm__30_,
  calc_stage_r_3__instr_operands__imm__29_,calc_stage_r_3__instr_operands__imm__28_,
  calc_stage_r_3__instr_operands__imm__27_,calc_stage_r_3__instr_operands__imm__26_,
  calc_stage_r_3__instr_operands__imm__25_,calc_stage_r_3__instr_operands__imm__24_,
  calc_stage_r_3__instr_operands__imm__23_,calc_stage_r_3__instr_operands__imm__22_,
  calc_stage_r_3__instr_operands__imm__21_,calc_stage_r_3__instr_operands__imm__20_,
  calc_stage_r_3__instr_operands__imm__19_,calc_stage_r_3__instr_operands__imm__18_,
  calc_stage_r_3__instr_operands__imm__17_,calc_stage_r_3__instr_operands__imm__16_,
  calc_stage_r_3__instr_operands__imm__15_,calc_stage_r_3__instr_operands__imm__14_,
  calc_stage_r_3__instr_operands__imm__13_,
  calc_stage_r_3__instr_operands__imm__12_,calc_stage_r_3__instr_operands__imm__11_,
  calc_stage_r_3__instr_operands__imm__10_,calc_stage_r_3__instr_operands__imm__9_,
  calc_stage_r_3__instr_operands__imm__8_,calc_stage_r_3__instr_operands__imm__7_,
  calc_stage_r_3__instr_operands__imm__6_,calc_stage_r_3__instr_operands__imm__5_,
  calc_stage_r_3__instr_operands__imm__4_,calc_stage_r_3__instr_operands__imm__3_,
  calc_stage_r_3__instr_operands__imm__2_,calc_stage_r_3__instr_operands__imm__1_,
  calc_stage_r_3__instr_operands__imm__0_,calc_stage_r_3__decode__instr_v_,calc_stage_r_3__decode__fe_nop_v_,
  calc_stage_r_3__decode__be_nop_v_,calc_stage_r_3__decode__me_nop_v_,
  calc_stage_r_3__decode__pipe_comp_v_,calc_stage_r_3__decode__pipe_int_v_,
  calc_stage_r_3__decode__pipe_mul_v_,calc_stage_r_3__decode__pipe_mem_v_,calc_stage_r_3__decode__pipe_fp_v_,
  calc_stage_r_3__decode__irf_w_v_,calc_stage_r_3__decode__frf_w_v_,
  calc_stage_r_3__decode__mhartid_r_v_,calc_stage_r_3__decode__dcache_w_v_,
  calc_stage_r_3__decode__dcache_r_v_,calc_stage_r_3__decode__fp_not_int_v_,
  calc_stage_r_3__decode__ret_v_,calc_stage_r_3__decode__amo_v_,calc_stage_r_3__decode__jmp_v_,
  calc_stage_r_3__decode__br_v_,calc_stage_r_3__decode__opw_v_,
  calc_stage_r_3__decode__fu_op__fu_op__3_,calc_stage_r_3__decode__fu_op__fu_op__2_,
  calc_stage_r_3__decode__fu_op__fu_op__1_,calc_stage_r_3__decode__fu_op__fu_op__0_,
  calc_stage_r_3__decode__rs1_addr__4_,calc_stage_r_3__decode__rs1_addr__3_,
  calc_stage_r_3__decode__rs1_addr__2_,calc_stage_r_3__decode__rs1_addr__1_,calc_stage_r_3__decode__rs1_addr__0_,
  calc_stage_r_3__decode__rs2_addr__4_,calc_stage_r_3__decode__rs2_addr__3_,
  calc_stage_r_3__decode__rs2_addr__2_,calc_stage_r_3__decode__rs2_addr__1_,
  calc_stage_r_3__decode__rs2_addr__0_,calc_stage_r_3__decode__src1_sel_,
  calc_stage_r_3__decode__src2_sel_,calc_stage_r_3__decode__baddr_sel_,calc_stage_r_3__decode__result_sel_,
  calc_stage_r_2__instr_metadata__itag__7_,
  calc_stage_r_2__instr_metadata__itag__6_,calc_stage_r_2__instr_metadata__itag__5_,
  calc_stage_r_2__instr_metadata__itag__4_,calc_stage_r_2__instr_metadata__itag__3_,
  calc_stage_r_2__instr_metadata__itag__2_,calc_stage_r_2__instr_metadata__itag__1_,
  calc_stage_r_2__instr_metadata__itag__0_,calc_stage_r_2__instr_metadata__fe_exception_not_instr_,
  calc_stage_r_2__instr_metadata__fe_exception_code__1_,
  calc_stage_r_2__instr_metadata__fe_exception_code__0_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__35_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__34_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__33_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__32_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__31_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__30_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__29_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__28_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__27_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__26_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__25_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__24_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__23_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__22_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__21_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__20_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__19_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__18_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__17_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__16_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__15_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__14_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__13_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__12_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__11_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__10_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__9_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__8_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__7_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__6_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__5_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__4_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__3_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__2_,calc_stage_r_2__instr_metadata__branch_metadata_fwd__1_,
  calc_stage_r_2__instr_metadata__branch_metadata_fwd__0_,calc_stage_r_2__instr__31_,
  calc_stage_r_2__instr__30_,calc_stage_r_2__instr__29_,
  calc_stage_r_2__instr__28_,calc_stage_r_2__instr__27_,calc_stage_r_2__instr__26_,
  calc_stage_r_2__instr__25_,calc_stage_r_2__instr__24_,calc_stage_r_2__instr__23_,
  calc_stage_r_2__instr__22_,calc_stage_r_2__instr__21_,calc_stage_r_2__instr__20_,
  calc_stage_r_2__instr__19_,calc_stage_r_2__instr__18_,calc_stage_r_2__instr__17_,
  calc_stage_r_2__instr__16_,calc_stage_r_2__instr__15_,calc_stage_r_2__instr__14_,
  calc_stage_r_2__instr__13_,calc_stage_r_2__instr__12_,calc_stage_r_2__instr__11_,
  calc_stage_r_2__instr__10_,calc_stage_r_2__instr__9_,calc_stage_r_2__instr__8_,
  calc_stage_r_2__instr__7_,calc_stage_r_2__instr__6_,calc_stage_r_2__instr__5_,
  calc_stage_r_2__instr__4_,calc_stage_r_2__instr__3_,calc_stage_r_2__instr__2_,
  calc_stage_r_2__instr__1_,calc_stage_r_2__instr__0_,calc_stage_r_2__instr_operands__rs1__63_,
  calc_stage_r_2__instr_operands__rs1__62_,calc_stage_r_2__instr_operands__rs1__61_,
  calc_stage_r_2__instr_operands__rs1__60_,calc_stage_r_2__instr_operands__rs1__59_,
  calc_stage_r_2__instr_operands__rs1__58_,calc_stage_r_2__instr_operands__rs1__57_,
  calc_stage_r_2__instr_operands__rs1__56_,calc_stage_r_2__instr_operands__rs1__55_,
  calc_stage_r_2__instr_operands__rs1__54_,calc_stage_r_2__instr_operands__rs1__53_,
  calc_stage_r_2__instr_operands__rs1__52_,calc_stage_r_2__instr_operands__rs1__51_,
  calc_stage_r_2__instr_operands__rs1__50_,
  calc_stage_r_2__instr_operands__rs1__49_,calc_stage_r_2__instr_operands__rs1__48_,
  calc_stage_r_2__instr_operands__rs1__47_,calc_stage_r_2__instr_operands__rs1__46_,
  calc_stage_r_2__instr_operands__rs1__45_,calc_stage_r_2__instr_operands__rs1__44_,
  calc_stage_r_2__instr_operands__rs1__43_,calc_stage_r_2__instr_operands__rs1__42_,
  calc_stage_r_2__instr_operands__rs1__41_,calc_stage_r_2__instr_operands__rs1__40_,
  calc_stage_r_2__instr_operands__rs1__39_,calc_stage_r_2__instr_operands__rs1__38_,
  calc_stage_r_2__instr_operands__rs1__37_,calc_stage_r_2__instr_operands__rs1__36_,
  calc_stage_r_2__instr_operands__rs1__35_,calc_stage_r_2__instr_operands__rs1__34_,
  calc_stage_r_2__instr_operands__rs1__33_,calc_stage_r_2__instr_operands__rs1__32_,
  calc_stage_r_2__instr_operands__rs1__31_,calc_stage_r_2__instr_operands__rs1__30_,
  calc_stage_r_2__instr_operands__rs1__29_,calc_stage_r_2__instr_operands__rs1__28_,
  calc_stage_r_2__instr_operands__rs1__27_,calc_stage_r_2__instr_operands__rs1__26_,
  calc_stage_r_2__instr_operands__rs1__25_,calc_stage_r_2__instr_operands__rs1__24_,
  calc_stage_r_2__instr_operands__rs1__23_,calc_stage_r_2__instr_operands__rs1__22_,
  calc_stage_r_2__instr_operands__rs1__21_,calc_stage_r_2__instr_operands__rs1__20_,
  calc_stage_r_2__instr_operands__rs1__19_,calc_stage_r_2__instr_operands__rs1__18_,
  calc_stage_r_2__instr_operands__rs1__17_,calc_stage_r_2__instr_operands__rs1__16_,
  calc_stage_r_2__instr_operands__rs1__15_,calc_stage_r_2__instr_operands__rs1__14_,
  calc_stage_r_2__instr_operands__rs1__13_,calc_stage_r_2__instr_operands__rs1__12_,
  calc_stage_r_2__instr_operands__rs1__11_,
  calc_stage_r_2__instr_operands__rs1__10_,calc_stage_r_2__instr_operands__rs1__9_,
  calc_stage_r_2__instr_operands__rs1__8_,calc_stage_r_2__instr_operands__rs1__7_,
  calc_stage_r_2__instr_operands__rs1__6_,calc_stage_r_2__instr_operands__rs1__5_,
  calc_stage_r_2__instr_operands__rs1__4_,calc_stage_r_2__instr_operands__rs1__3_,
  calc_stage_r_2__instr_operands__rs1__2_,calc_stage_r_2__instr_operands__rs1__1_,
  calc_stage_r_2__instr_operands__rs1__0_,calc_stage_r_2__instr_operands__rs2__63_,
  calc_stage_r_2__instr_operands__rs2__62_,calc_stage_r_2__instr_operands__rs2__61_,
  calc_stage_r_2__instr_operands__rs2__60_,calc_stage_r_2__instr_operands__rs2__59_,
  calc_stage_r_2__instr_operands__rs2__58_,calc_stage_r_2__instr_operands__rs2__57_,
  calc_stage_r_2__instr_operands__rs2__56_,calc_stage_r_2__instr_operands__rs2__55_,
  calc_stage_r_2__instr_operands__rs2__54_,calc_stage_r_2__instr_operands__rs2__53_,
  calc_stage_r_2__instr_operands__rs2__52_,calc_stage_r_2__instr_operands__rs2__51_,
  calc_stage_r_2__instr_operands__rs2__50_,calc_stage_r_2__instr_operands__rs2__49_,
  calc_stage_r_2__instr_operands__rs2__48_,calc_stage_r_2__instr_operands__rs2__47_,
  calc_stage_r_2__instr_operands__rs2__46_,calc_stage_r_2__instr_operands__rs2__45_,
  calc_stage_r_2__instr_operands__rs2__44_,calc_stage_r_2__instr_operands__rs2__43_,
  calc_stage_r_2__instr_operands__rs2__42_,calc_stage_r_2__instr_operands__rs2__41_,
  calc_stage_r_2__instr_operands__rs2__40_,calc_stage_r_2__instr_operands__rs2__39_,
  calc_stage_r_2__instr_operands__rs2__38_,calc_stage_r_2__instr_operands__rs2__37_,
  calc_stage_r_2__instr_operands__rs2__36_,calc_stage_r_2__instr_operands__rs2__35_,
  calc_stage_r_2__instr_operands__rs2__34_,calc_stage_r_2__instr_operands__rs2__33_,
  calc_stage_r_2__instr_operands__rs2__32_,calc_stage_r_2__instr_operands__rs2__31_,
  calc_stage_r_2__instr_operands__rs2__30_,calc_stage_r_2__instr_operands__rs2__29_,
  calc_stage_r_2__instr_operands__rs2__28_,calc_stage_r_2__instr_operands__rs2__27_,
  calc_stage_r_2__instr_operands__rs2__26_,calc_stage_r_2__instr_operands__rs2__25_,
  calc_stage_r_2__instr_operands__rs2__24_,
  calc_stage_r_2__instr_operands__rs2__23_,calc_stage_r_2__instr_operands__rs2__22_,
  calc_stage_r_2__instr_operands__rs2__21_,calc_stage_r_2__instr_operands__rs2__20_,
  calc_stage_r_2__instr_operands__rs2__19_,calc_stage_r_2__instr_operands__rs2__18_,
  calc_stage_r_2__instr_operands__rs2__17_,calc_stage_r_2__instr_operands__rs2__16_,
  calc_stage_r_2__instr_operands__rs2__15_,calc_stage_r_2__instr_operands__rs2__14_,
  calc_stage_r_2__instr_operands__rs2__13_,calc_stage_r_2__instr_operands__rs2__12_,
  calc_stage_r_2__instr_operands__rs2__11_,calc_stage_r_2__instr_operands__rs2__10_,
  calc_stage_r_2__instr_operands__rs2__9_,calc_stage_r_2__instr_operands__rs2__8_,
  calc_stage_r_2__instr_operands__rs2__7_,calc_stage_r_2__instr_operands__rs2__6_,
  calc_stage_r_2__instr_operands__rs2__5_,calc_stage_r_2__instr_operands__rs2__4_,
  calc_stage_r_2__instr_operands__rs2__3_,exc_stage_r_3__poison_v_,exc_stage_r_3__roll_v_,
  exc_stage_r_3__illegal_instr_v_,exc_stage_r_3__tlb_miss_v_,exc_stage_r_3__load_fault_v_,
  exc_stage_r_3__store_fault_v_,exc_stage_r_3__cache_miss_v_,exc_stage_r_2__poison_v_,
  exc_stage_r_2__roll_v_,exc_stage_r_2__illegal_instr_v_,exc_stage_r_2__tlb_miss_v_,
  exc_stage_r_2__load_fault_v_,exc_stage_r_2__store_fault_v_,
  exc_stage_r_2__cache_miss_v_,exc_stage_r_1__poison_v_,exc_stage_r_1__roll_v_,
  exc_stage_r_1__illegal_instr_v_,exc_stage_r_1__tlb_miss_v_,exc_stage_r_1__load_fault_v_,
  exc_stage_r_1__store_fault_v_,exc_stage_r_1__cache_miss_v_,exc_stage_r_0__poison_v_,
  exc_stage_r_0__roll_v_,exc_stage_r_0__illegal_instr_v_,exc_stage_r_0__tlb_miss_v_,
  exc_stage_r_0__load_fault_v_,exc_stage_r_0__store_fault_v_,exc_stage_r_0__cache_miss_v_,
  n_7_net_,n_14_net_,n_15_net_,issue_pkt_r_instr__31_,issue_pkt_r_instr__30_,
  issue_pkt_r_instr__29_,issue_pkt_r_instr__28_,issue_pkt_r_instr__27_,
  issue_pkt_r_instr__26_,issue_pkt_r_instr__25_,issue_pkt_r_instr__24_,issue_pkt_r_instr__23_,
  issue_pkt_r_instr__22_,issue_pkt_r_instr__21_,issue_pkt_r_instr__20_,
  issue_pkt_r_instr__19_,issue_pkt_r_instr__18_,issue_pkt_r_instr__17_,issue_pkt_r_instr__16_,
  issue_pkt_r_instr__15_,issue_pkt_r_instr__14_,issue_pkt_r_instr__13_,
  issue_pkt_r_instr__12_,issue_pkt_r_instr__11_,issue_pkt_r_instr__10_,issue_pkt_r_instr__9_,
  issue_pkt_r_instr__8_,issue_pkt_r_instr__7_,issue_pkt_r_instr__6_,issue_pkt_r_instr__5_,
  issue_pkt_r_instr__4_,issue_pkt_r_instr__3_,issue_pkt_r_instr__2_,
  issue_pkt_r_instr__1_,issue_pkt_r_instr__0_,n_16_net_,n_17_net_,n_18_net_,n_19_net_,n_20_net_,
  int_calc_result_result__63_,int_calc_result_result__62_,
  int_calc_result_result__61_,int_calc_result_result__60_,int_calc_result_result__59_,
  int_calc_result_result__58_,int_calc_result_result__57_,int_calc_result_result__56_,
  int_calc_result_result__55_,int_calc_result_result__54_,int_calc_result_result__53_,
  int_calc_result_result__52_,int_calc_result_result__51_,int_calc_result_result__50_,
  int_calc_result_result__49_,int_calc_result_result__48_,int_calc_result_result__47_,
  int_calc_result_result__46_,int_calc_result_result__45_,int_calc_result_result__44_,
  int_calc_result_result__43_,int_calc_result_result__42_,
  int_calc_result_result__41_,int_calc_result_result__40_,int_calc_result_result__39_,
  int_calc_result_result__38_,int_calc_result_result__37_,int_calc_result_result__36_,
  int_calc_result_result__35_,int_calc_result_result__34_,int_calc_result_result__33_,
  int_calc_result_result__32_,int_calc_result_result__31_,int_calc_result_result__30_,
  int_calc_result_result__29_,int_calc_result_result__28_,int_calc_result_result__27_,
  int_calc_result_result__26_,int_calc_result_result__25_,int_calc_result_result__24_,
  int_calc_result_result__23_,int_calc_result_result__22_,
  int_calc_result_result__21_,int_calc_result_result__20_,int_calc_result_result__19_,
  int_calc_result_result__18_,int_calc_result_result__17_,int_calc_result_result__16_,
  int_calc_result_result__15_,int_calc_result_result__14_,int_calc_result_result__13_,
  int_calc_result_result__12_,int_calc_result_result__11_,int_calc_result_result__10_,
  int_calc_result_result__9_,int_calc_result_result__8_,int_calc_result_result__7_,
  int_calc_result_result__6_,int_calc_result_result__5_,int_calc_result_result__4_,
  int_calc_result_result__3_,int_calc_result_result__2_,int_calc_result_result__1_,
  int_calc_result_result__0_,calc_stage_r_2__instr_operands__rs2__2_,
  calc_stage_r_2__instr_operands__rs2__1_,calc_stage_r_2__instr_operands__rs2__0_,
  calc_stage_r_2__instr_operands__imm__63_,calc_stage_r_2__instr_operands__imm__62_,
  calc_stage_r_2__instr_operands__imm__61_,calc_stage_r_2__instr_operands__imm__60_,
  calc_stage_r_2__instr_operands__imm__59_,calc_stage_r_2__instr_operands__imm__58_,
  calc_stage_r_2__instr_operands__imm__57_,calc_stage_r_2__instr_operands__imm__56_,
  calc_stage_r_2__instr_operands__imm__55_,calc_stage_r_2__instr_operands__imm__54_,
  calc_stage_r_2__instr_operands__imm__53_,calc_stage_r_2__instr_operands__imm__52_,
  calc_stage_r_2__instr_operands__imm__51_,calc_stage_r_2__instr_operands__imm__50_,
  calc_stage_r_2__instr_operands__imm__49_,calc_stage_r_2__instr_operands__imm__48_,
  calc_stage_r_2__instr_operands__imm__47_,calc_stage_r_2__instr_operands__imm__46_,
  calc_stage_r_2__instr_operands__imm__45_,
  calc_stage_r_2__instr_operands__imm__44_,calc_stage_r_2__instr_operands__imm__43_,
  calc_stage_r_2__instr_operands__imm__42_,calc_stage_r_2__instr_operands__imm__41_,
  calc_stage_r_2__instr_operands__imm__40_,calc_stage_r_2__instr_operands__imm__39_,
  calc_stage_r_2__instr_operands__imm__38_,calc_stage_r_2__instr_operands__imm__37_,
  calc_stage_r_2__instr_operands__imm__36_,calc_stage_r_2__instr_operands__imm__35_,
  calc_stage_r_2__instr_operands__imm__34_,calc_stage_r_2__instr_operands__imm__33_,
  calc_stage_r_2__instr_operands__imm__32_,calc_stage_r_2__instr_operands__imm__31_,
  calc_stage_r_2__instr_operands__imm__30_,calc_stage_r_2__instr_operands__imm__29_,
  calc_stage_r_2__instr_operands__imm__28_,calc_stage_r_2__instr_operands__imm__27_,
  calc_stage_r_2__instr_operands__imm__26_,calc_stage_r_2__instr_operands__imm__25_,
  calc_stage_r_2__instr_operands__imm__24_,calc_stage_r_2__instr_operands__imm__23_,
  calc_stage_r_2__instr_operands__imm__22_,calc_stage_r_2__instr_operands__imm__21_,
  calc_stage_r_2__instr_operands__imm__20_,calc_stage_r_2__instr_operands__imm__19_,
  calc_stage_r_2__instr_operands__imm__18_,calc_stage_r_2__instr_operands__imm__17_,
  calc_stage_r_2__instr_operands__imm__16_,calc_stage_r_2__instr_operands__imm__15_,
  calc_stage_r_2__instr_operands__imm__14_,calc_stage_r_2__instr_operands__imm__13_,
  calc_stage_r_2__instr_operands__imm__12_,calc_stage_r_2__instr_operands__imm__11_,
  calc_stage_r_2__instr_operands__imm__10_,calc_stage_r_2__instr_operands__imm__9_,
  calc_stage_r_2__instr_operands__imm__8_,calc_stage_r_2__instr_operands__imm__7_,
  calc_stage_r_2__instr_operands__imm__6_,calc_stage_r_2__instr_operands__imm__5_,
  calc_stage_r_2__instr_operands__imm__4_,calc_stage_r_2__instr_operands__imm__3_,
  calc_stage_r_2__instr_operands__imm__2_,calc_stage_r_2__instr_operands__imm__1_,
  calc_stage_r_2__instr_operands__imm__0_,calc_stage_r_2__decode__instr_v_,
  calc_stage_r_2__decode__fe_nop_v_,calc_stage_r_2__decode__be_nop_v_,
  calc_stage_r_2__decode__me_nop_v_,calc_stage_r_2__decode__pipe_comp_v_,
  calc_stage_r_2__decode__pipe_int_v_,calc_stage_r_2__decode__pipe_mul_v_,calc_stage_r_2__decode__pipe_mem_v_,
  calc_stage_r_2__decode__pipe_fp_v_,calc_stage_r_2__decode__irf_w_v_,
  calc_stage_r_2__decode__frf_w_v_,calc_stage_r_2__decode__mhartid_r_v_,
  calc_stage_r_2__decode__dcache_w_v_,calc_stage_r_2__decode__dcache_r_v_,
  calc_stage_r_2__decode__fp_not_int_v_,calc_stage_r_2__decode__amo_v_,calc_stage_r_2__decode__jmp_v_,
  calc_stage_r_2__decode__br_v_,calc_stage_r_2__decode__opw_v_,
  calc_stage_r_2__decode__fu_op__fu_op__3_,calc_stage_r_2__decode__fu_op__fu_op__2_,
  calc_stage_r_2__decode__fu_op__fu_op__1_,calc_stage_r_2__decode__fu_op__fu_op__0_,
  calc_stage_r_2__decode__rs1_addr__4_,calc_stage_r_2__decode__rs1_addr__3_,
  calc_stage_r_2__decode__rs1_addr__2_,calc_stage_r_2__decode__rs1_addr__1_,calc_stage_r_2__decode__rs1_addr__0_,
  calc_stage_r_2__decode__rs2_addr__4_,calc_stage_r_2__decode__rs2_addr__3_,
  calc_stage_r_2__decode__rs2_addr__2_,calc_stage_r_2__decode__rs2_addr__1_,
  calc_stage_r_2__decode__rs2_addr__0_,calc_stage_r_2__decode__src1_sel_,
  calc_stage_r_2__decode__src2_sel_,calc_stage_r_2__decode__baddr_sel_,calc_stage_r_2__decode__result_sel_,
  calc_stage_r_1__instr_metadata__itag__7_,
  calc_stage_r_1__instr_metadata__itag__6_,calc_stage_r_1__instr_metadata__itag__5_,
  calc_stage_r_1__instr_metadata__itag__4_,calc_stage_r_1__instr_metadata__itag__3_,
  calc_stage_r_1__instr_metadata__itag__2_,calc_stage_r_1__instr_metadata__itag__1_,
  calc_stage_r_1__instr_metadata__itag__0_,calc_stage_r_1__instr_metadata__pc__63_,
  calc_stage_r_1__instr_metadata__pc__62_,calc_stage_r_1__instr_metadata__pc__61_,
  calc_stage_r_1__instr_metadata__pc__60_,calc_stage_r_1__instr_metadata__pc__59_,
  calc_stage_r_1__instr_metadata__pc__58_,calc_stage_r_1__instr_metadata__pc__57_,
  calc_stage_r_1__instr_metadata__pc__56_,calc_stage_r_1__instr_metadata__pc__55_,
  calc_stage_r_1__instr_metadata__pc__54_,calc_stage_r_1__instr_metadata__pc__53_,
  calc_stage_r_1__instr_metadata__pc__52_,calc_stage_r_1__instr_metadata__pc__51_,
  calc_stage_r_1__instr_metadata__pc__50_,calc_stage_r_1__instr_metadata__pc__49_,
  calc_stage_r_1__instr_metadata__pc__48_,calc_stage_r_1__instr_metadata__pc__47_,
  calc_stage_r_1__instr_metadata__pc__46_,calc_stage_r_1__instr_metadata__pc__45_,
  calc_stage_r_1__instr_metadata__pc__44_,calc_stage_r_1__instr_metadata__pc__43_,
  calc_stage_r_1__instr_metadata__pc__42_,calc_stage_r_1__instr_metadata__pc__41_,
  calc_stage_r_1__instr_metadata__pc__40_,calc_stage_r_1__instr_metadata__pc__39_,
  calc_stage_r_1__instr_metadata__pc__38_,calc_stage_r_1__instr_metadata__pc__37_,
  calc_stage_r_1__instr_metadata__pc__36_,calc_stage_r_1__instr_metadata__pc__35_,
  calc_stage_r_1__instr_metadata__pc__34_,calc_stage_r_1__instr_metadata__pc__33_,
  calc_stage_r_1__instr_metadata__pc__32_,calc_stage_r_1__instr_metadata__pc__31_,
  calc_stage_r_1__instr_metadata__pc__30_,calc_stage_r_1__instr_metadata__pc__29_,
  calc_stage_r_1__instr_metadata__pc__28_,calc_stage_r_1__instr_metadata__pc__27_,
  calc_stage_r_1__instr_metadata__pc__26_,calc_stage_r_1__instr_metadata__pc__25_,
  calc_stage_r_1__instr_metadata__pc__24_,calc_stage_r_1__instr_metadata__pc__23_,
  calc_stage_r_1__instr_metadata__pc__22_,calc_stage_r_1__instr_metadata__pc__21_,
  calc_stage_r_1__instr_metadata__pc__20_,calc_stage_r_1__instr_metadata__pc__19_,
  calc_stage_r_1__instr_metadata__pc__18_,calc_stage_r_1__instr_metadata__pc__17_,
  calc_stage_r_1__instr_metadata__pc__16_,calc_stage_r_1__instr_metadata__pc__15_,
  calc_stage_r_1__instr_metadata__pc__14_,calc_stage_r_1__instr_metadata__pc__13_,
  calc_stage_r_1__instr_metadata__pc__12_,calc_stage_r_1__instr_metadata__pc__11_,
  calc_stage_r_1__instr_metadata__pc__10_,calc_stage_r_1__instr_metadata__pc__9_,
  calc_stage_r_1__instr_metadata__pc__8_,calc_stage_r_1__instr_metadata__pc__7_,
  calc_stage_r_1__instr_metadata__pc__6_,calc_stage_r_1__instr_metadata__pc__5_,
  calc_stage_r_1__instr_metadata__pc__4_,calc_stage_r_1__instr_metadata__pc__3_,calc_stage_r_1__instr_metadata__pc__2_,
  calc_stage_r_1__instr_metadata__pc__1_,calc_stage_r_1__instr_metadata__pc__0_,
  calc_stage_r_1__instr_metadata__fe_exception_not_instr_,
  calc_stage_r_1__instr_metadata__fe_exception_code__1_,
  calc_stage_r_1__instr_metadata__fe_exception_code__0_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__35_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__34_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__33_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__32_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__31_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__30_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__29_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__28_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__27_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__26_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__25_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__24_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__23_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__22_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__21_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__20_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__19_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__18_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__17_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__16_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__15_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__14_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__13_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__12_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__11_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__10_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__9_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__8_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__7_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__6_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__5_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__4_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__3_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__2_,calc_stage_r_1__instr_metadata__branch_metadata_fwd__1_,
  calc_stage_r_1__instr_metadata__branch_metadata_fwd__0_,calc_stage_r_1__instr__31_,
  calc_stage_r_1__instr__30_,calc_stage_r_1__instr__29_,calc_stage_r_1__instr__28_,
  calc_stage_r_1__instr__27_,calc_stage_r_1__instr__26_,calc_stage_r_1__instr__25_,
  calc_stage_r_1__instr__24_,calc_stage_r_1__instr__23_,calc_stage_r_1__instr__22_,
  calc_stage_r_1__instr__21_,calc_stage_r_1__instr__20_,calc_stage_r_1__instr__19_,
  calc_stage_r_1__instr__18_,calc_stage_r_1__instr__17_,calc_stage_r_1__instr__16_,
  calc_stage_r_1__instr__15_,calc_stage_r_1__instr__14_,calc_stage_r_1__instr__13_,
  calc_stage_r_1__instr__12_,calc_stage_r_1__instr__11_,calc_stage_r_1__instr__10_,
  calc_stage_r_1__instr__9_,calc_stage_r_1__instr__8_,calc_stage_r_1__instr__7_,
  calc_stage_r_1__instr__6_,calc_stage_r_1__instr__5_,calc_stage_r_1__instr__4_,
  calc_stage_r_1__instr__3_,calc_stage_r_1__instr__2_,calc_stage_r_1__instr__1_,
  calc_stage_r_1__instr__0_,calc_stage_r_1__instr_operands__rs1__63_,
  calc_stage_r_1__instr_operands__rs1__62_,calc_stage_r_1__instr_operands__rs1__61_,
  calc_stage_r_1__instr_operands__rs1__60_,calc_stage_r_1__instr_operands__rs1__59_,
  calc_stage_r_1__instr_operands__rs1__58_,calc_stage_r_1__instr_operands__rs1__57_,
  calc_stage_r_1__instr_operands__rs1__56_,calc_stage_r_1__instr_operands__rs1__55_,
  calc_stage_r_1__instr_operands__rs1__54_,calc_stage_r_1__instr_operands__rs1__53_,
  calc_stage_r_1__instr_operands__rs1__52_,calc_stage_r_1__instr_operands__rs1__51_,
  calc_stage_r_1__instr_operands__rs1__50_,calc_stage_r_1__instr_operands__rs1__49_,
  calc_stage_r_1__instr_operands__rs1__48_,calc_stage_r_1__instr_operands__rs1__47_,
  calc_stage_r_1__instr_operands__rs1__46_,calc_stage_r_1__instr_operands__rs1__45_,
  calc_stage_r_1__instr_operands__rs1__44_,calc_stage_r_1__instr_operands__rs1__43_,
  calc_stage_r_1__instr_operands__rs1__42_,
  calc_stage_r_1__instr_operands__rs1__41_,calc_stage_r_1__instr_operands__rs1__40_,
  calc_stage_r_1__instr_operands__rs1__39_,calc_stage_r_1__instr_operands__rs1__38_,
  calc_stage_r_1__instr_operands__rs1__37_,calc_stage_r_1__instr_operands__rs1__36_,
  calc_stage_r_1__instr_operands__rs1__35_,calc_stage_r_1__instr_operands__rs1__34_,
  calc_stage_r_1__instr_operands__rs1__33_,calc_stage_r_1__instr_operands__rs1__32_,
  calc_stage_r_1__instr_operands__rs1__31_,calc_stage_r_1__instr_operands__rs1__30_,
  calc_stage_r_1__instr_operands__rs1__29_,calc_stage_r_1__instr_operands__rs1__28_,
  calc_stage_r_1__instr_operands__rs1__27_,calc_stage_r_1__instr_operands__rs1__26_,
  calc_stage_r_1__instr_operands__rs1__25_,calc_stage_r_1__instr_operands__rs1__24_,
  calc_stage_r_1__instr_operands__rs1__23_,calc_stage_r_1__instr_operands__rs1__22_,
  calc_stage_r_1__instr_operands__rs1__21_,calc_stage_r_1__instr_operands__rs1__20_,
  calc_stage_r_1__instr_operands__rs1__19_,calc_stage_r_1__instr_operands__rs1__18_,
  calc_stage_r_1__instr_operands__rs1__17_,calc_stage_r_1__instr_operands__rs1__16_,
  calc_stage_r_1__instr_operands__rs1__15_,calc_stage_r_1__instr_operands__rs1__14_,
  calc_stage_r_1__instr_operands__rs1__13_,calc_stage_r_1__instr_operands__rs1__12_,
  calc_stage_r_1__instr_operands__rs1__11_,calc_stage_r_1__instr_operands__rs1__10_,
  calc_stage_r_1__instr_operands__rs1__9_,calc_stage_r_1__instr_operands__rs1__8_,
  calc_stage_r_1__instr_operands__rs1__7_,calc_stage_r_1__instr_operands__rs1__6_,
  calc_stage_r_1__instr_operands__rs1__5_,calc_stage_r_1__instr_operands__rs1__4_,
  calc_stage_r_1__instr_operands__rs1__3_,calc_stage_r_1__instr_operands__rs1__2_,
  calc_stage_r_1__instr_operands__rs1__1_,calc_stage_r_1__instr_operands__rs1__0_,
  calc_stage_r_1__instr_operands__rs2__63_,calc_stage_r_1__instr_operands__rs2__62_,
  calc_stage_r_1__instr_operands__rs2__61_,calc_stage_r_1__instr_operands__rs2__60_,
  calc_stage_r_1__instr_operands__rs2__59_,calc_stage_r_1__instr_operands__rs2__58_,
  calc_stage_r_1__instr_operands__rs2__57_,calc_stage_r_1__instr_operands__rs2__56_,
  calc_stage_r_1__instr_operands__rs2__55_,
  calc_stage_r_1__instr_operands__rs2__54_,calc_stage_r_1__instr_operands__rs2__53_,
  calc_stage_r_1__instr_operands__rs2__52_,calc_stage_r_1__instr_operands__rs2__51_,
  calc_stage_r_1__instr_operands__rs2__50_,calc_stage_r_1__instr_operands__rs2__49_,
  calc_stage_r_1__instr_operands__rs2__48_,calc_stage_r_1__instr_operands__rs2__47_,
  calc_stage_r_1__instr_operands__rs2__46_,calc_stage_r_1__instr_operands__rs2__45_,
  calc_stage_r_1__instr_operands__rs2__44_,calc_stage_r_1__instr_operands__rs2__43_,
  calc_stage_r_1__instr_operands__rs2__42_,calc_stage_r_1__instr_operands__rs2__41_,
  calc_stage_r_1__instr_operands__rs2__40_,calc_stage_r_1__instr_operands__rs2__39_,
  calc_stage_r_1__instr_operands__rs2__38_,calc_stage_r_1__instr_operands__rs2__37_,
  calc_stage_r_1__instr_operands__rs2__36_,calc_stage_r_1__instr_operands__rs2__35_,
  calc_stage_r_1__instr_operands__rs2__34_,calc_stage_r_1__instr_operands__rs2__33_,
  calc_stage_r_1__instr_operands__rs2__32_,calc_stage_r_1__instr_operands__rs2__31_,
  calc_stage_r_1__instr_operands__rs2__30_,calc_stage_r_1__instr_operands__rs2__29_,
  calc_stage_r_1__instr_operands__rs2__28_,calc_stage_r_1__instr_operands__rs2__27_,
  calc_stage_r_1__instr_operands__rs2__26_,calc_stage_r_1__instr_operands__rs2__25_,
  calc_stage_r_1__instr_operands__rs2__24_,calc_stage_r_1__instr_operands__rs2__23_,
  calc_stage_r_1__instr_operands__rs2__22_,calc_stage_r_1__instr_operands__rs2__21_,
  calc_stage_r_1__instr_operands__rs2__20_,calc_stage_r_1__instr_operands__rs2__19_,
  calc_stage_r_1__instr_operands__rs2__18_,calc_stage_r_1__instr_operands__rs2__17_,
  calc_stage_r_1__instr_operands__rs2__16_,
  calc_stage_r_1__instr_operands__rs2__15_,calc_stage_r_1__instr_operands__rs2__14_,
  calc_stage_r_1__instr_operands__rs2__13_,calc_stage_r_1__instr_operands__rs2__12_,
  calc_stage_r_1__instr_operands__rs2__11_,calc_stage_r_1__instr_operands__rs2__10_,
  calc_stage_r_1__instr_operands__rs2__9_,calc_stage_r_1__instr_operands__rs2__8_,
  calc_stage_r_1__instr_operands__rs2__7_,calc_stage_r_1__instr_operands__rs2__6_,
  calc_stage_r_1__instr_operands__rs2__5_,calc_stage_r_1__instr_operands__rs2__4_,
  calc_stage_r_1__instr_operands__rs2__3_,calc_stage_r_1__instr_operands__rs2__2_,
  calc_stage_r_1__instr_operands__rs2__1_,calc_stage_r_1__instr_operands__rs2__0_,
  calc_stage_r_1__instr_operands__imm__63_,calc_stage_r_1__instr_operands__imm__62_,
  calc_stage_r_1__instr_operands__imm__61_,calc_stage_r_1__instr_operands__imm__60_,
  calc_stage_r_1__instr_operands__imm__59_,calc_stage_r_1__instr_operands__imm__58_,
  calc_stage_r_1__instr_operands__imm__57_,calc_stage_r_1__instr_operands__imm__56_,
  calc_stage_r_1__instr_operands__imm__55_,calc_stage_r_1__instr_operands__imm__54_,
  calc_stage_r_1__instr_operands__imm__53_,calc_stage_r_1__instr_operands__imm__52_,
  calc_stage_r_1__instr_operands__imm__51_,calc_stage_r_1__instr_operands__imm__50_,
  calc_stage_r_1__instr_operands__imm__49_,calc_stage_r_1__instr_operands__imm__48_,
  calc_stage_r_1__instr_operands__imm__47_,calc_stage_r_1__instr_operands__imm__46_,
  calc_stage_r_1__instr_operands__imm__45_,calc_stage_r_1__instr_operands__imm__44_,
  calc_stage_r_1__instr_operands__imm__43_,calc_stage_r_1__instr_operands__imm__42_,
  calc_stage_r_1__instr_operands__imm__41_,calc_stage_r_1__instr_operands__imm__40_,
  calc_stage_r_1__instr_operands__imm__39_,calc_stage_r_1__instr_operands__imm__38_,
  calc_stage_r_1__instr_operands__imm__37_,calc_stage_r_1__instr_operands__imm__36_,
  calc_stage_r_1__instr_operands__imm__35_,calc_stage_r_1__instr_operands__imm__34_,
  calc_stage_r_1__instr_operands__imm__33_,calc_stage_r_1__instr_operands__imm__32_,
  calc_stage_r_1__instr_operands__imm__31_,calc_stage_r_1__instr_operands__imm__30_,
  calc_stage_r_1__instr_operands__imm__29_,
  calc_stage_r_1__instr_operands__imm__28_,calc_stage_r_1__instr_operands__imm__27_,
  calc_stage_r_1__instr_operands__imm__26_,calc_stage_r_1__instr_operands__imm__25_,
  calc_stage_r_1__instr_operands__imm__24_,calc_stage_r_1__instr_operands__imm__23_,
  calc_stage_r_1__instr_operands__imm__22_,calc_stage_r_1__instr_operands__imm__21_,
  calc_stage_r_1__instr_operands__imm__20_,calc_stage_r_1__instr_operands__imm__19_,
  calc_stage_r_1__instr_operands__imm__18_,calc_stage_r_1__instr_operands__imm__17_,
  calc_stage_r_1__instr_operands__imm__16_,calc_stage_r_1__instr_operands__imm__15_,
  calc_stage_r_1__instr_operands__imm__14_,calc_stage_r_1__instr_operands__imm__13_,
  calc_stage_r_1__instr_operands__imm__12_,calc_stage_r_1__instr_operands__imm__11_,
  calc_stage_r_1__instr_operands__imm__10_,calc_stage_r_1__instr_operands__imm__9_,
  calc_stage_r_1__instr_operands__imm__8_,calc_stage_r_1__instr_operands__imm__7_,
  calc_stage_r_1__instr_operands__imm__6_,calc_stage_r_1__instr_operands__imm__5_,
  calc_stage_r_1__instr_operands__imm__4_,calc_stage_r_1__instr_operands__imm__3_,
  calc_stage_r_1__instr_operands__imm__2_,calc_stage_r_1__instr_operands__imm__1_,
  calc_stage_r_1__instr_operands__imm__0_,calc_stage_r_1__decode__instr_v_,
  calc_stage_r_1__decode__fe_nop_v_,calc_stage_r_1__decode__be_nop_v_,calc_stage_r_1__decode__me_nop_v_,
  calc_stage_r_1__decode__pipe_comp_v_,calc_stage_r_1__decode__pipe_int_v_,
  calc_stage_r_1__decode__pipe_mul_v_,calc_stage_r_1__decode__pipe_mem_v_,
  calc_stage_r_1__decode__pipe_fp_v_,calc_stage_r_1__decode__irf_w_v_,
  calc_stage_r_1__decode__frf_w_v_,calc_stage_r_1__decode__mhartid_r_v_,calc_stage_r_1__decode__dcache_w_v_,
  calc_stage_r_1__decode__dcache_r_v_,calc_stage_r_1__decode__fp_not_int_v_,
  calc_stage_r_1__decode__ret_v_,calc_stage_r_1__decode__amo_v_,
  calc_stage_r_1__decode__jmp_v_,calc_stage_r_1__decode__br_v_,calc_stage_r_1__decode__opw_v_,
  calc_stage_r_1__decode__fu_op__fu_op__3_,calc_stage_r_1__decode__fu_op__fu_op__2_,
  calc_stage_r_1__decode__fu_op__fu_op__1_,calc_stage_r_1__decode__fu_op__fu_op__0_,
  calc_stage_r_1__decode__rs1_addr__4_,calc_stage_r_1__decode__rs1_addr__3_,
  calc_stage_r_1__decode__rs1_addr__2_,calc_stage_r_1__decode__rs1_addr__1_,
  calc_stage_r_1__decode__rs1_addr__0_,calc_stage_r_1__decode__rs2_addr__4_,
  calc_stage_r_1__decode__rs2_addr__3_,calc_stage_r_1__decode__rs2_addr__2_,calc_stage_r_1__decode__rs2_addr__1_,
  calc_stage_r_1__decode__rs2_addr__0_,calc_stage_r_1__decode__src1_sel_,
  calc_stage_r_1__decode__src2_sel_,calc_stage_r_1__decode__baddr_sel_,
  calc_stage_r_1__decode__result_sel_,calc_stage_r_0__instr_metadata__itag__7_,
  calc_stage_r_0__instr_metadata__itag__6_,calc_stage_r_0__instr_metadata__itag__5_,
  calc_stage_r_0__instr_metadata__itag__4_,calc_stage_r_0__instr_metadata__itag__3_,
  calc_stage_r_0__instr_metadata__itag__2_,calc_stage_r_0__instr_metadata__itag__1_,
  calc_stage_r_0__instr_metadata__itag__0_,calc_stage_r_0__instr_metadata__pc__63_,
  calc_stage_r_0__instr_metadata__pc__62_,calc_stage_r_0__instr_metadata__pc__61_,
  calc_stage_r_0__instr_metadata__pc__60_,calc_stage_r_0__instr_metadata__pc__59_,
  calc_stage_r_0__instr_metadata__pc__58_,calc_stage_r_0__instr_metadata__pc__57_,
  calc_stage_r_0__instr_metadata__pc__56_,calc_stage_r_0__instr_metadata__pc__55_,
  calc_stage_r_0__instr_metadata__pc__54_,calc_stage_r_0__instr_metadata__pc__53_,
  calc_stage_r_0__instr_metadata__pc__52_,calc_stage_r_0__instr_metadata__pc__51_,
  calc_stage_r_0__instr_metadata__pc__50_,calc_stage_r_0__instr_metadata__pc__49_,
  calc_stage_r_0__instr_metadata__pc__48_,calc_stage_r_0__instr_metadata__pc__47_,
  calc_stage_r_0__instr_metadata__pc__46_,calc_stage_r_0__instr_metadata__pc__45_,
  calc_stage_r_0__instr_metadata__pc__44_,calc_stage_r_0__instr_metadata__pc__43_,
  calc_stage_r_0__instr_metadata__pc__42_,calc_stage_r_0__instr_metadata__pc__41_,
  calc_stage_r_0__instr_metadata__pc__40_,calc_stage_r_0__instr_metadata__pc__39_,
  calc_stage_r_0__instr_metadata__pc__38_,calc_stage_r_0__instr_metadata__pc__37_,
  calc_stage_r_0__instr_metadata__pc__36_,calc_stage_r_0__instr_metadata__pc__35_,
  calc_stage_r_0__instr_metadata__pc__34_,calc_stage_r_0__instr_metadata__pc__33_,
  calc_stage_r_0__instr_metadata__pc__32_,calc_stage_r_0__instr_metadata__pc__31_,
  calc_stage_r_0__instr_metadata__pc__30_,calc_stage_r_0__instr_metadata__pc__29_,
  calc_stage_r_0__instr_metadata__pc__28_,calc_stage_r_0__instr_metadata__pc__27_,
  calc_stage_r_0__instr_metadata__pc__26_,calc_stage_r_0__instr_metadata__pc__25_,
  calc_stage_r_0__instr_metadata__pc__24_,calc_stage_r_0__instr_metadata__pc__23_,
  calc_stage_r_0__instr_metadata__pc__22_,calc_stage_r_0__instr_metadata__pc__21_,
  calc_stage_r_0__instr_metadata__pc__20_,calc_stage_r_0__instr_metadata__pc__19_,
  calc_stage_r_0__instr_metadata__pc__18_,calc_stage_r_0__instr_metadata__pc__17_,
  calc_stage_r_0__instr_metadata__pc__16_,calc_stage_r_0__instr_metadata__pc__15_,
  calc_stage_r_0__instr_metadata__pc__14_,calc_stage_r_0__instr_metadata__pc__13_,
  calc_stage_r_0__instr_metadata__pc__12_,calc_stage_r_0__instr_metadata__pc__11_,
  calc_stage_r_0__instr_metadata__pc__10_,calc_stage_r_0__instr_metadata__pc__9_,
  calc_stage_r_0__instr_metadata__pc__8_,calc_stage_r_0__instr_metadata__pc__7_,
  calc_stage_r_0__instr_metadata__pc__6_,calc_stage_r_0__instr_metadata__pc__5_,
  calc_stage_r_0__instr_metadata__pc__4_,calc_stage_r_0__instr_metadata__pc__3_,
  calc_stage_r_0__instr_metadata__pc__2_,calc_stage_r_0__instr_metadata__pc__1_,
  calc_stage_r_0__instr_metadata__pc__0_,calc_stage_r_0__instr_metadata__fe_exception_not_instr_,
  calc_stage_r_0__instr_metadata__fe_exception_code__1_,
  calc_stage_r_0__instr_metadata__fe_exception_code__0_,calc_stage_r_0__instr__31_,calc_stage_r_0__instr__30_,
  calc_stage_r_0__instr__29_,calc_stage_r_0__instr__28_,calc_stage_r_0__instr__27_,
  calc_stage_r_0__instr__26_,calc_stage_r_0__instr__25_,calc_stage_r_0__instr__24_,
  calc_stage_r_0__instr__23_,calc_stage_r_0__instr__22_,calc_stage_r_0__instr__21_,
  calc_stage_r_0__instr__20_,calc_stage_r_0__instr__19_,calc_stage_r_0__instr__18_,
  calc_stage_r_0__instr__17_,calc_stage_r_0__instr__16_,calc_stage_r_0__instr__15_,
  calc_stage_r_0__instr__14_,calc_stage_r_0__instr__13_,calc_stage_r_0__instr__12_,
  calc_stage_r_0__instr__11_,calc_stage_r_0__instr__10_,calc_stage_r_0__instr__9_,
  calc_stage_r_0__instr__8_,calc_stage_r_0__instr__7_,calc_stage_r_0__instr__6_,
  calc_stage_r_0__instr__5_,calc_stage_r_0__instr__4_,calc_stage_r_0__instr__3_,
  calc_stage_r_0__instr__2_,calc_stage_r_0__instr__1_,calc_stage_r_0__instr__0_,
  calc_stage_r_0__instr_operands__rs1__63_,calc_stage_r_0__instr_operands__rs1__62_,
  calc_stage_r_0__instr_operands__rs1__61_,calc_stage_r_0__instr_operands__rs1__60_,
  calc_stage_r_0__instr_operands__rs1__59_,calc_stage_r_0__instr_operands__rs1__58_,
  calc_stage_r_0__instr_operands__rs1__57_,calc_stage_r_0__instr_operands__rs1__56_,
  calc_stage_r_0__instr_operands__rs1__55_,
  calc_stage_r_0__instr_operands__rs1__54_,calc_stage_r_0__instr_operands__rs1__53_,
  calc_stage_r_0__instr_operands__rs1__52_,calc_stage_r_0__instr_operands__rs1__51_,
  calc_stage_r_0__instr_operands__rs1__50_,calc_stage_r_0__instr_operands__rs1__49_,
  calc_stage_r_0__instr_operands__rs1__48_,calc_stage_r_0__instr_operands__rs1__47_,
  calc_stage_r_0__instr_operands__rs1__46_,calc_stage_r_0__instr_operands__rs1__45_,
  calc_stage_r_0__instr_operands__rs1__44_,calc_stage_r_0__instr_operands__rs1__43_,
  calc_stage_r_0__instr_operands__rs1__42_,calc_stage_r_0__instr_operands__rs1__41_,
  calc_stage_r_0__instr_operands__rs1__40_,calc_stage_r_0__instr_operands__rs1__39_,
  calc_stage_r_0__instr_operands__rs1__38_,calc_stage_r_0__instr_operands__rs1__37_,
  calc_stage_r_0__instr_operands__rs1__36_,calc_stage_r_0__instr_operands__rs1__35_,
  calc_stage_r_0__instr_operands__rs1__34_,calc_stage_r_0__instr_operands__rs1__33_,
  calc_stage_r_0__instr_operands__rs1__32_,calc_stage_r_0__instr_operands__rs1__31_,
  calc_stage_r_0__instr_operands__rs1__30_,calc_stage_r_0__instr_operands__rs1__29_,
  calc_stage_r_0__instr_operands__rs1__28_,calc_stage_r_0__instr_operands__rs1__27_,
  calc_stage_r_0__instr_operands__rs1__26_,calc_stage_r_0__instr_operands__rs1__25_,
  calc_stage_r_0__instr_operands__rs1__24_,calc_stage_r_0__instr_operands__rs1__23_,
  calc_stage_r_0__instr_operands__rs1__22_,calc_stage_r_0__instr_operands__rs1__21_,
  calc_stage_r_0__instr_operands__rs1__20_,calc_stage_r_0__instr_operands__rs1__19_,
  calc_stage_r_0__instr_operands__rs1__18_,calc_stage_r_0__instr_operands__rs1__17_,
  calc_stage_r_0__instr_operands__rs1__16_,calc_stage_r_0__instr_operands__rs1__15_,
  calc_stage_r_0__instr_operands__rs1__14_,
  calc_stage_r_0__instr_operands__rs1__13_,calc_stage_r_0__instr_operands__rs1__12_,
  calc_stage_r_0__instr_operands__rs1__11_,calc_stage_r_0__instr_operands__rs1__10_,
  calc_stage_r_0__instr_operands__rs1__9_,calc_stage_r_0__instr_operands__rs1__8_,
  calc_stage_r_0__instr_operands__rs1__7_,calc_stage_r_0__instr_operands__rs1__6_,
  calc_stage_r_0__instr_operands__rs1__5_,calc_stage_r_0__instr_operands__rs1__4_,
  calc_stage_r_0__instr_operands__rs1__3_,calc_stage_r_0__instr_operands__rs1__2_,
  calc_stage_r_0__instr_operands__rs1__1_,calc_stage_r_0__instr_operands__rs1__0_,
  calc_stage_r_0__instr_operands__rs2__63_,calc_stage_r_0__instr_operands__rs2__62_,
  calc_stage_r_0__instr_operands__rs2__61_,calc_stage_r_0__instr_operands__rs2__60_,
  calc_stage_r_0__instr_operands__rs2__59_,calc_stage_r_0__instr_operands__rs2__58_,
  calc_stage_r_0__instr_operands__rs2__57_,calc_stage_r_0__instr_operands__rs2__56_,
  calc_stage_r_0__instr_operands__rs2__55_,calc_stage_r_0__instr_operands__rs2__54_,
  calc_stage_r_0__instr_operands__rs2__53_,calc_stage_r_0__instr_operands__rs2__52_,
  calc_stage_r_0__instr_operands__rs2__51_,calc_stage_r_0__instr_operands__rs2__50_,
  calc_stage_r_0__instr_operands__rs2__49_,calc_stage_r_0__instr_operands__rs2__48_,
  calc_stage_r_0__instr_operands__rs2__47_,calc_stage_r_0__instr_operands__rs2__46_,
  calc_stage_r_0__instr_operands__rs2__45_,calc_stage_r_0__instr_operands__rs2__44_,
  calc_stage_r_0__instr_operands__rs2__43_,calc_stage_r_0__instr_operands__rs2__42_,
  calc_stage_r_0__instr_operands__rs2__41_,calc_stage_r_0__instr_operands__rs2__40_,
  calc_stage_r_0__instr_operands__rs2__39_,calc_stage_r_0__instr_operands__rs2__38_,
  calc_stage_r_0__instr_operands__rs2__37_,calc_stage_r_0__instr_operands__rs2__36_,
  calc_stage_r_0__instr_operands__rs2__35_,calc_stage_r_0__instr_operands__rs2__34_,
  calc_stage_r_0__instr_operands__rs2__33_,calc_stage_r_0__instr_operands__rs2__32_,
  calc_stage_r_0__instr_operands__rs2__31_,calc_stage_r_0__instr_operands__rs2__30_,
  calc_stage_r_0__instr_operands__rs2__29_,
  calc_stage_r_0__instr_operands__rs2__28_,calc_stage_r_0__instr_operands__rs2__27_,
  calc_stage_r_0__instr_operands__rs2__26_,calc_stage_r_0__instr_operands__rs2__25_,
  calc_stage_r_0__instr_operands__rs2__24_,calc_stage_r_0__instr_operands__rs2__23_,
  calc_stage_r_0__instr_operands__rs2__22_,calc_stage_r_0__instr_operands__rs2__21_,
  calc_stage_r_0__instr_operands__rs2__20_,calc_stage_r_0__instr_operands__rs2__19_,
  calc_stage_r_0__instr_operands__rs2__18_,calc_stage_r_0__instr_operands__rs2__17_,
  calc_stage_r_0__instr_operands__rs2__16_,calc_stage_r_0__instr_operands__rs2__15_,
  calc_stage_r_0__instr_operands__rs2__14_,calc_stage_r_0__instr_operands__rs2__13_,
  calc_stage_r_0__instr_operands__rs2__12_,calc_stage_r_0__instr_operands__rs2__11_,
  calc_stage_r_0__instr_operands__rs2__10_,calc_stage_r_0__instr_operands__rs2__9_,
  calc_stage_r_0__instr_operands__rs2__8_,calc_stage_r_0__instr_operands__rs2__7_,
  calc_stage_r_0__instr_operands__rs2__6_,calc_stage_r_0__instr_operands__rs2__5_,
  calc_stage_r_0__instr_operands__rs2__4_,calc_stage_r_0__instr_operands__rs2__3_,
  calc_stage_r_0__instr_operands__rs2__2_,calc_stage_r_0__instr_operands__rs2__1_,
  calc_stage_r_0__instr_operands__rs2__0_,calc_stage_r_0__instr_operands__imm__63_,
  calc_stage_r_0__instr_operands__imm__62_,calc_stage_r_0__instr_operands__imm__61_,
  calc_stage_r_0__instr_operands__imm__60_,calc_stage_r_0__instr_operands__imm__59_,
  calc_stage_r_0__instr_operands__imm__58_,calc_stage_r_0__instr_operands__imm__57_,
  calc_stage_r_0__instr_operands__imm__56_,calc_stage_r_0__instr_operands__imm__55_,
  calc_stage_r_0__instr_operands__imm__54_,calc_stage_r_0__instr_operands__imm__53_,
  calc_stage_r_0__instr_operands__imm__52_,calc_stage_r_0__instr_operands__imm__51_,
  calc_stage_r_0__instr_operands__imm__50_,calc_stage_r_0__instr_operands__imm__49_,
  calc_stage_r_0__instr_operands__imm__48_,calc_stage_r_0__instr_operands__imm__47_,
  calc_stage_r_0__instr_operands__imm__46_,calc_stage_r_0__instr_operands__imm__45_,
  calc_stage_r_0__instr_operands__imm__44_,calc_stage_r_0__instr_operands__imm__43_,
  calc_stage_r_0__instr_operands__imm__42_,
  calc_stage_r_0__instr_operands__imm__41_,calc_stage_r_0__instr_operands__imm__40_,
  calc_stage_r_0__instr_operands__imm__39_,calc_stage_r_0__instr_operands__imm__38_,
  calc_stage_r_0__instr_operands__imm__37_,calc_stage_r_0__instr_operands__imm__36_,
  calc_stage_r_0__instr_operands__imm__35_,calc_stage_r_0__instr_operands__imm__34_,
  calc_stage_r_0__instr_operands__imm__33_,calc_stage_r_0__instr_operands__imm__32_,
  calc_stage_r_0__instr_operands__imm__31_,calc_stage_r_0__instr_operands__imm__30_,
  calc_stage_r_0__instr_operands__imm__29_,calc_stage_r_0__instr_operands__imm__28_,
  calc_stage_r_0__instr_operands__imm__27_,calc_stage_r_0__instr_operands__imm__26_,
  calc_stage_r_0__instr_operands__imm__25_,calc_stage_r_0__instr_operands__imm__24_,
  calc_stage_r_0__instr_operands__imm__23_,calc_stage_r_0__instr_operands__imm__22_,
  calc_stage_r_0__instr_operands__imm__21_,calc_stage_r_0__instr_operands__imm__20_,
  calc_stage_r_0__instr_operands__imm__19_,calc_stage_r_0__instr_operands__imm__18_,
  calc_stage_r_0__instr_operands__imm__17_,calc_stage_r_0__instr_operands__imm__16_,
  calc_stage_r_0__instr_operands__imm__15_,calc_stage_r_0__instr_operands__imm__14_,
  calc_stage_r_0__instr_operands__imm__13_,calc_stage_r_0__instr_operands__imm__12_,
  calc_stage_r_0__instr_operands__imm__11_,calc_stage_r_0__instr_operands__imm__10_,
  calc_stage_r_0__instr_operands__imm__9_,calc_stage_r_0__instr_operands__imm__8_,
  calc_stage_r_0__instr_operands__imm__7_,calc_stage_r_0__instr_operands__imm__6_,
  calc_stage_r_0__instr_operands__imm__5_,calc_stage_r_0__instr_operands__imm__4_,
  calc_stage_r_0__instr_operands__imm__3_,calc_stage_r_0__instr_operands__imm__2_,
  calc_stage_r_0__instr_operands__imm__1_,calc_stage_r_0__instr_operands__imm__0_,
  calc_stage_r_0__decode__instr_v_,calc_stage_r_0__decode__fe_nop_v_,
  calc_stage_r_0__decode__be_nop_v_,calc_stage_r_0__decode__me_nop_v_,
  calc_stage_r_0__decode__pipe_comp_v_,calc_stage_r_0__decode__pipe_int_v_,calc_stage_r_0__decode__pipe_mul_v_,
  calc_stage_r_0__decode__pipe_mem_v_,calc_stage_r_0__decode__pipe_fp_v_,
  calc_stage_r_0__decode__irf_w_v_,calc_stage_r_0__decode__frf_w_v_,
  calc_stage_r_0__decode__mhartid_r_v_,calc_stage_r_0__decode__dcache_w_v_,
  calc_stage_r_0__decode__dcache_r_v_,calc_stage_r_0__decode__fp_not_int_v_,calc_stage_r_0__decode__ret_v_,
  calc_stage_r_0__decode__amo_v_,calc_stage_r_0__decode__jmp_v_,
  calc_stage_r_0__decode__br_v_,calc_stage_r_0__decode__opw_v_,calc_stage_r_0__decode__fu_op__fu_op__3_,
  calc_stage_r_0__decode__fu_op__fu_op__2_,calc_stage_r_0__decode__fu_op__fu_op__1_,
  calc_stage_r_0__decode__fu_op__fu_op__0_,calc_stage_r_0__decode__rs1_addr__4_,
  calc_stage_r_0__decode__rs1_addr__3_,calc_stage_r_0__decode__rs1_addr__2_,
  calc_stage_r_0__decode__rs1_addr__1_,calc_stage_r_0__decode__rs1_addr__0_,
  calc_stage_r_0__decode__rs2_addr__4_,calc_stage_r_0__decode__rs2_addr__3_,
  calc_stage_r_0__decode__rs2_addr__2_,calc_stage_r_0__decode__rs2_addr__1_,
  calc_stage_r_0__decode__rs2_addr__0_,calc_stage_r_0__decode__src1_sel_,calc_stage_r_0__decode__src2_sel_,
  calc_stage_r_0__decode__baddr_sel_,calc_stage_r_0__decode__result_sel_,
  dispatch_pkt_instr_metadata__itag__7_,dispatch_pkt_instr_metadata__itag__6_,
  dispatch_pkt_instr_metadata__itag__5_,dispatch_pkt_instr_metadata__itag__4_,
  dispatch_pkt_instr_metadata__itag__3_,dispatch_pkt_instr_metadata__itag__2_,
  dispatch_pkt_instr_metadata__itag__1_,dispatch_pkt_instr_metadata__itag__0_,
  dispatch_pkt_instr_metadata__fe_exception_not_instr_,dispatch_pkt_instr_metadata__fe_exception_code__1_,
  dispatch_pkt_instr_metadata__fe_exception_code__0_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__35_,dispatch_pkt_instr_metadata__branch_metadata_fwd__34_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__33_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__32_,dispatch_pkt_instr_metadata__branch_metadata_fwd__31_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__30_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__29_,dispatch_pkt_instr_metadata__branch_metadata_fwd__28_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__27_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__26_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__25_,dispatch_pkt_instr_metadata__branch_metadata_fwd__24_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__23_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__22_,dispatch_pkt_instr_metadata__branch_metadata_fwd__21_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__20_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__19_,dispatch_pkt_instr_metadata__branch_metadata_fwd__18_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__17_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__16_,dispatch_pkt_instr_metadata__branch_metadata_fwd__15_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__14_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__13_,dispatch_pkt_instr_metadata__branch_metadata_fwd__12_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__11_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__10_,dispatch_pkt_instr_metadata__branch_metadata_fwd__9_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__8_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__7_,dispatch_pkt_instr_metadata__branch_metadata_fwd__6_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__5_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__4_,dispatch_pkt_instr_metadata__branch_metadata_fwd__3_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__2_,
  dispatch_pkt_instr_metadata__branch_metadata_fwd__1_,dispatch_pkt_instr_metadata__branch_metadata_fwd__0_,
  dispatch_pkt_instr_operands__rs1__63_,dispatch_pkt_instr_operands__rs1__62_,
  dispatch_pkt_instr_operands__rs1__61_,dispatch_pkt_instr_operands__rs1__60_,
  dispatch_pkt_instr_operands__rs1__59_,dispatch_pkt_instr_operands__rs1__58_,
  dispatch_pkt_instr_operands__rs1__57_,dispatch_pkt_instr_operands__rs1__56_,
  dispatch_pkt_instr_operands__rs1__55_,dispatch_pkt_instr_operands__rs1__54_,dispatch_pkt_instr_operands__rs1__53_,
  dispatch_pkt_instr_operands__rs1__52_,dispatch_pkt_instr_operands__rs1__51_,
  dispatch_pkt_instr_operands__rs1__50_,dispatch_pkt_instr_operands__rs1__49_,
  dispatch_pkt_instr_operands__rs1__48_,dispatch_pkt_instr_operands__rs1__47_,
  dispatch_pkt_instr_operands__rs1__46_,dispatch_pkt_instr_operands__rs1__45_,
  dispatch_pkt_instr_operands__rs1__44_,dispatch_pkt_instr_operands__rs1__43_,
  dispatch_pkt_instr_operands__rs1__42_,dispatch_pkt_instr_operands__rs1__41_,
  dispatch_pkt_instr_operands__rs1__40_,dispatch_pkt_instr_operands__rs1__39_,
  dispatch_pkt_instr_operands__rs1__38_,dispatch_pkt_instr_operands__rs1__37_,
  dispatch_pkt_instr_operands__rs1__36_,dispatch_pkt_instr_operands__rs1__35_,
  dispatch_pkt_instr_operands__rs1__34_,dispatch_pkt_instr_operands__rs1__33_,dispatch_pkt_instr_operands__rs1__32_,
  dispatch_pkt_instr_operands__rs1__31_,dispatch_pkt_instr_operands__rs1__30_,
  dispatch_pkt_instr_operands__rs1__29_,dispatch_pkt_instr_operands__rs1__28_,
  dispatch_pkt_instr_operands__rs1__27_,dispatch_pkt_instr_operands__rs1__26_,
  dispatch_pkt_instr_operands__rs1__25_,dispatch_pkt_instr_operands__rs1__24_,
  dispatch_pkt_instr_operands__rs1__23_,dispatch_pkt_instr_operands__rs1__22_,
  dispatch_pkt_instr_operands__rs1__21_,dispatch_pkt_instr_operands__rs1__20_,
  dispatch_pkt_instr_operands__rs1__19_,dispatch_pkt_instr_operands__rs1__18_,
  dispatch_pkt_instr_operands__rs1__17_,dispatch_pkt_instr_operands__rs1__16_,
  dispatch_pkt_instr_operands__rs1__15_,dispatch_pkt_instr_operands__rs1__14_,dispatch_pkt_instr_operands__rs1__13_,
  dispatch_pkt_instr_operands__rs1__12_,dispatch_pkt_instr_operands__rs1__11_,
  dispatch_pkt_instr_operands__rs1__10_,dispatch_pkt_instr_operands__rs1__9_,
  dispatch_pkt_instr_operands__rs1__8_,dispatch_pkt_instr_operands__rs1__7_,
  dispatch_pkt_instr_operands__rs1__6_,dispatch_pkt_instr_operands__rs1__5_,
  dispatch_pkt_instr_operands__rs1__4_,dispatch_pkt_instr_operands__rs1__3_,
  dispatch_pkt_instr_operands__rs1__2_,dispatch_pkt_instr_operands__rs1__1_,
  dispatch_pkt_instr_operands__rs1__0_,dispatch_pkt_instr_operands__rs2__63_,dispatch_pkt_instr_operands__rs2__62_,
  dispatch_pkt_instr_operands__rs2__61_,dispatch_pkt_instr_operands__rs2__60_,
  dispatch_pkt_instr_operands__rs2__59_,dispatch_pkt_instr_operands__rs2__58_,
  dispatch_pkt_instr_operands__rs2__57_,dispatch_pkt_instr_operands__rs2__56_,
  dispatch_pkt_instr_operands__rs2__55_,dispatch_pkt_instr_operands__rs2__54_,
  dispatch_pkt_instr_operands__rs2__53_,dispatch_pkt_instr_operands__rs2__52_,
  dispatch_pkt_instr_operands__rs2__51_,dispatch_pkt_instr_operands__rs2__50_,
  dispatch_pkt_instr_operands__rs2__49_,dispatch_pkt_instr_operands__rs2__48_,
  dispatch_pkt_instr_operands__rs2__47_,dispatch_pkt_instr_operands__rs2__46_,
  dispatch_pkt_instr_operands__rs2__45_,dispatch_pkt_instr_operands__rs2__44_,
  dispatch_pkt_instr_operands__rs2__43_,dispatch_pkt_instr_operands__rs2__42_,dispatch_pkt_instr_operands__rs2__41_,
  dispatch_pkt_instr_operands__rs2__40_,dispatch_pkt_instr_operands__rs2__39_,
  dispatch_pkt_instr_operands__rs2__38_,dispatch_pkt_instr_operands__rs2__37_,
  dispatch_pkt_instr_operands__rs2__36_,dispatch_pkt_instr_operands__rs2__35_,
  dispatch_pkt_instr_operands__rs2__34_,dispatch_pkt_instr_operands__rs2__33_,
  dispatch_pkt_instr_operands__rs2__32_,dispatch_pkt_instr_operands__rs2__31_,
  dispatch_pkt_instr_operands__rs2__30_,dispatch_pkt_instr_operands__rs2__29_,
  dispatch_pkt_instr_operands__rs2__28_,dispatch_pkt_instr_operands__rs2__27_,
  dispatch_pkt_instr_operands__rs2__26_,dispatch_pkt_instr_operands__rs2__25_,
  dispatch_pkt_instr_operands__rs2__24_,dispatch_pkt_instr_operands__rs2__23_,dispatch_pkt_instr_operands__rs2__22_,
  dispatch_pkt_instr_operands__rs2__21_,dispatch_pkt_instr_operands__rs2__20_,
  dispatch_pkt_instr_operands__rs2__19_,dispatch_pkt_instr_operands__rs2__18_,
  dispatch_pkt_instr_operands__rs2__17_,dispatch_pkt_instr_operands__rs2__16_,
  dispatch_pkt_instr_operands__rs2__15_,dispatch_pkt_instr_operands__rs2__14_,
  dispatch_pkt_instr_operands__rs2__13_,dispatch_pkt_instr_operands__rs2__12_,
  dispatch_pkt_instr_operands__rs2__11_,dispatch_pkt_instr_operands__rs2__10_,
  dispatch_pkt_instr_operands__rs2__9_,dispatch_pkt_instr_operands__rs2__8_,
  dispatch_pkt_instr_operands__rs2__7_,dispatch_pkt_instr_operands__rs2__6_,dispatch_pkt_instr_operands__rs2__5_,
  dispatch_pkt_instr_operands__rs2__4_,dispatch_pkt_instr_operands__rs2__3_,
  dispatch_pkt_instr_operands__rs2__2_,dispatch_pkt_instr_operands__rs2__1_,
  dispatch_pkt_instr_operands__rs2__0_,dispatch_pkt_instr_operands__imm__63_,
  dispatch_pkt_instr_operands__imm__62_,dispatch_pkt_instr_operands__imm__61_,
  dispatch_pkt_instr_operands__imm__60_,dispatch_pkt_instr_operands__imm__59_,
  dispatch_pkt_instr_operands__imm__58_,dispatch_pkt_instr_operands__imm__57_,
  dispatch_pkt_instr_operands__imm__56_,dispatch_pkt_instr_operands__imm__55_,
  dispatch_pkt_instr_operands__imm__54_,dispatch_pkt_instr_operands__imm__53_,
  dispatch_pkt_instr_operands__imm__52_,dispatch_pkt_instr_operands__imm__51_,dispatch_pkt_instr_operands__imm__50_,
  dispatch_pkt_instr_operands__imm__49_,dispatch_pkt_instr_operands__imm__48_,
  dispatch_pkt_instr_operands__imm__47_,dispatch_pkt_instr_operands__imm__46_,
  dispatch_pkt_instr_operands__imm__45_,dispatch_pkt_instr_operands__imm__44_,
  dispatch_pkt_instr_operands__imm__43_,dispatch_pkt_instr_operands__imm__42_,
  dispatch_pkt_instr_operands__imm__41_,dispatch_pkt_instr_operands__imm__40_,
  dispatch_pkt_instr_operands__imm__39_,dispatch_pkt_instr_operands__imm__38_,
  dispatch_pkt_instr_operands__imm__37_,dispatch_pkt_instr_operands__imm__36_,
  dispatch_pkt_instr_operands__imm__35_,dispatch_pkt_instr_operands__imm__34_,
  dispatch_pkt_instr_operands__imm__33_,dispatch_pkt_instr_operands__imm__32_,dispatch_pkt_instr_operands__imm__31_,
  dispatch_pkt_instr_operands__imm__30_,dispatch_pkt_instr_operands__imm__29_,
  dispatch_pkt_instr_operands__imm__28_,dispatch_pkt_instr_operands__imm__27_,
  dispatch_pkt_instr_operands__imm__26_,dispatch_pkt_instr_operands__imm__25_,
  dispatch_pkt_instr_operands__imm__24_,dispatch_pkt_instr_operands__imm__23_,
  dispatch_pkt_instr_operands__imm__22_,dispatch_pkt_instr_operands__imm__21_,
  dispatch_pkt_instr_operands__imm__20_,dispatch_pkt_instr_operands__imm__19_,
  dispatch_pkt_instr_operands__imm__18_,dispatch_pkt_instr_operands__imm__17_,
  dispatch_pkt_instr_operands__imm__16_,dispatch_pkt_instr_operands__imm__15_,
  dispatch_pkt_instr_operands__imm__14_,dispatch_pkt_instr_operands__imm__13_,
  dispatch_pkt_instr_operands__imm__12_,dispatch_pkt_instr_operands__imm__11_,dispatch_pkt_instr_operands__imm__10_,
  dispatch_pkt_instr_operands__imm__9_,dispatch_pkt_instr_operands__imm__8_,
  dispatch_pkt_instr_operands__imm__7_,dispatch_pkt_instr_operands__imm__6_,
  dispatch_pkt_instr_operands__imm__5_,dispatch_pkt_instr_operands__imm__4_,
  dispatch_pkt_instr_operands__imm__3_,dispatch_pkt_instr_operands__imm__2_,
  dispatch_pkt_instr_operands__imm__1_,dispatch_pkt_instr_operands__imm__0_,dispatch_pkt_decode__instr_v_,
  dispatch_pkt_decode__fe_nop_v_,dispatch_pkt_decode__be_nop_v_,
  dispatch_pkt_decode__me_nop_v_,dispatch_pkt_decode__pipe_comp_v_,dispatch_pkt_decode__pipe_int_v_,
  dispatch_pkt_decode__pipe_mul_v_,dispatch_pkt_decode__pipe_mem_v_,
  dispatch_pkt_decode__pipe_fp_v_,dispatch_pkt_decode__irf_w_v_,dispatch_pkt_decode__frf_w_v_,
  dispatch_pkt_decode__mhartid_r_v_,dispatch_pkt_decode__dcache_w_v_,
  dispatch_pkt_decode__dcache_r_v_,dispatch_pkt_decode__ret_v_,dispatch_pkt_decode__amo_v_,
  dispatch_pkt_decode__jmp_v_,dispatch_pkt_decode__br_v_,dispatch_pkt_decode__opw_v_,
  dispatch_pkt_decode__rd_addr__4_,dispatch_pkt_decode__rd_addr__3_,
  dispatch_pkt_decode__rd_addr__2_,dispatch_pkt_decode__rd_addr__1_,dispatch_pkt_decode__rd_addr__0_,
  dispatch_pkt_decode__src1_sel_,dispatch_pkt_decode__src2_sel_,
  dispatch_pkt_decode__baddr_sel_,dispatch_pkt_decode__result_sel_,exc_stage_n_3__roll_v_,
  exc_stage_n_3__cache_miss_v_,exc_stage_n_2__poison_v_,exc_stage_n_2__roll_v_,
  exc_stage_n_1__poison_v_,exc_stage_n_1__roll_v_,exc_stage_n_0__illegal_instr_v_,N0,N1,N2,N3,
  N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,
  N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,
  N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,
  N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,
  N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,
  N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,
  N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,
  N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,
  N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,
  N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,
  N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,
  N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,
  N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,
  N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,
  N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
  N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,
  N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309;
  wire [63:0] irf_rs1,irf_rs2,frf_rs1,frf_rs2,bypass_irs1,bypass_irs2,bypass_frs1,bypass_frs2;
  wire [4:1] comp_stage_n_slice_iwb_v,comp_stage_n_slice_fwb_v;
  wire [639:0] comp_stage_n;
  assign calc_status_o[2] = 1'b0;
  assign cmt_trace_stage_reg_o[8] = calc_status_o[113];
  assign cmt_trace_stage_reg_o[7] = calc_status_o[112];
  assign cmt_trace_stage_reg_o[6] = calc_status_o[111];
  assign cmt_trace_stage_reg_o[5] = calc_status_o[110];
  assign cmt_trace_stage_reg_o[4] = calc_status_o[109];

  bp_be_regfile
  int_regfile
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .issue_v_i(issue_pkt_v_i),
    .dispatch_v_i(chk_dispatch_v_i),
    .rd_w_v_i(n_0_net_),
    .rd_addr_i(calc_status_o[103:99]),
    .rd_data_i({ comp_stage_r_3__result__63_, comp_stage_r_3__result__62_, comp_stage_r_3__result__61_, comp_stage_r_3__result__60_, comp_stage_r_3__result__59_, comp_stage_r_3__result__58_, comp_stage_r_3__result__57_, comp_stage_r_3__result__56_, comp_stage_r_3__result__55_, comp_stage_r_3__result__54_, comp_stage_r_3__result__53_, comp_stage_r_3__result__52_, comp_stage_r_3__result__51_, comp_stage_r_3__result__50_, comp_stage_r_3__result__49_, comp_stage_r_3__result__48_, comp_stage_r_3__result__47_, comp_stage_r_3__result__46_, comp_stage_r_3__result__45_, comp_stage_r_3__result__44_, comp_stage_r_3__result__43_, comp_stage_r_3__result__42_, comp_stage_r_3__result__41_, comp_stage_r_3__result__40_, comp_stage_r_3__result__39_, comp_stage_r_3__result__38_, comp_stage_r_3__result__37_, comp_stage_r_3__result__36_, comp_stage_r_3__result__35_, comp_stage_r_3__result__34_, comp_stage_r_3__result__33_, comp_stage_r_3__result__32_, comp_stage_r_3__result__31_, comp_stage_r_3__result__30_, comp_stage_r_3__result__29_, comp_stage_r_3__result__28_, comp_stage_r_3__result__27_, comp_stage_r_3__result__26_, comp_stage_r_3__result__25_, comp_stage_r_3__result__24_, comp_stage_r_3__result__23_, comp_stage_r_3__result__22_, comp_stage_r_3__result__21_, comp_stage_r_3__result__20_, comp_stage_r_3__result__19_, comp_stage_r_3__result__18_, comp_stage_r_3__result__17_, comp_stage_r_3__result__16_, comp_stage_r_3__result__15_, comp_stage_r_3__result__14_, comp_stage_r_3__result__13_, comp_stage_r_3__result__12_, comp_stage_r_3__result__11_, comp_stage_r_3__result__10_, comp_stage_r_3__result__9_, comp_stage_r_3__result__8_, comp_stage_r_3__result__7_, comp_stage_r_3__result__6_, comp_stage_r_3__result__5_, comp_stage_r_3__result__4_, comp_stage_r_3__result__3_, comp_stage_r_3__result__2_, comp_stage_r_3__result__1_, comp_stage_r_3__result__0_ }),
    .rs1_r_v_i(issue_pkt_i[77]),
    .rs1_addr_i(issue_pkt_i[73:69]),
    .rs1_data_o(irf_rs1),
    .rs2_r_v_i(issue_pkt_i[76]),
    .rs2_addr_i(issue_pkt_i[68:64]),
    .rs2_data_o(irf_rs2)
  );


  bp_be_regfile
  float_regfile
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .issue_v_i(issue_pkt_v_i),
    .dispatch_v_i(chk_dispatch_v_i),
    .rd_w_v_i(n_7_net_),
    .rd_addr_i(calc_status_o[113:109]),
    .rd_data_i(cmt_trace_result_o[127:64]),
    .rs1_r_v_i(issue_pkt_i[75]),
    .rs1_addr_i(issue_pkt_i[73:69]),
    .rs1_data_o(frf_rs1),
    .rs2_r_v_i(issue_pkt_i[74]),
    .rs2_addr_i(issue_pkt_i[68:64]),
    .rs2_data_o(frf_rs2)
  );


  bsg_dff_reset_en_width_p221
  issue_reg
  (
    .clk_i(clk_i),
    .reset_i(n_14_net_),
    .en_i(n_15_net_),
    .data_i(issue_pkt_i),
    .data_o({ dispatch_pkt_instr_metadata__itag__7_, dispatch_pkt_instr_metadata__itag__6_, dispatch_pkt_instr_metadata__itag__5_, dispatch_pkt_instr_metadata__itag__4_, dispatch_pkt_instr_metadata__itag__3_, dispatch_pkt_instr_metadata__itag__2_, dispatch_pkt_instr_metadata__itag__1_, dispatch_pkt_instr_metadata__itag__0_, calc_status_o[300:237], dispatch_pkt_instr_metadata__fe_exception_not_instr_, dispatch_pkt_instr_metadata__fe_exception_code__1_, dispatch_pkt_instr_metadata__fe_exception_code__0_, dispatch_pkt_instr_metadata__branch_metadata_fwd__35_, dispatch_pkt_instr_metadata__branch_metadata_fwd__34_, dispatch_pkt_instr_metadata__branch_metadata_fwd__33_, dispatch_pkt_instr_metadata__branch_metadata_fwd__32_, dispatch_pkt_instr_metadata__branch_metadata_fwd__31_, dispatch_pkt_instr_metadata__branch_metadata_fwd__30_, dispatch_pkt_instr_metadata__branch_metadata_fwd__29_, dispatch_pkt_instr_metadata__branch_metadata_fwd__28_, dispatch_pkt_instr_metadata__branch_metadata_fwd__27_, dispatch_pkt_instr_metadata__branch_metadata_fwd__26_, dispatch_pkt_instr_metadata__branch_metadata_fwd__25_, dispatch_pkt_instr_metadata__branch_metadata_fwd__24_, dispatch_pkt_instr_metadata__branch_metadata_fwd__23_, dispatch_pkt_instr_metadata__branch_metadata_fwd__22_, dispatch_pkt_instr_metadata__branch_metadata_fwd__21_, dispatch_pkt_instr_metadata__branch_metadata_fwd__20_, dispatch_pkt_instr_metadata__branch_metadata_fwd__19_, dispatch_pkt_instr_metadata__branch_metadata_fwd__18_, dispatch_pkt_instr_metadata__branch_metadata_fwd__17_, dispatch_pkt_instr_metadata__branch_metadata_fwd__16_, dispatch_pkt_instr_metadata__branch_metadata_fwd__15_, dispatch_pkt_instr_metadata__branch_metadata_fwd__14_, dispatch_pkt_instr_metadata__branch_metadata_fwd__13_, dispatch_pkt_instr_metadata__branch_metadata_fwd__12_, dispatch_pkt_instr_metadata__branch_metadata_fwd__11_, dispatch_pkt_instr_metadata__branch_metadata_fwd__10_, dispatch_pkt_instr_metadata__branch_metadata_fwd__9_, dispatch_pkt_instr_metadata__branch_metadata_fwd__8_, dispatch_pkt_instr_metadata__branch_metadata_fwd__7_, dispatch_pkt_instr_metadata__branch_metadata_fwd__6_, dispatch_pkt_instr_metadata__branch_metadata_fwd__5_, dispatch_pkt_instr_metadata__branch_metadata_fwd__4_, dispatch_pkt_instr_metadata__branch_metadata_fwd__3_, dispatch_pkt_instr_metadata__branch_metadata_fwd__2_, dispatch_pkt_instr_metadata__branch_metadata_fwd__1_, dispatch_pkt_instr_metadata__branch_metadata_fwd__0_, issue_pkt_r_instr__31_, issue_pkt_r_instr__30_, issue_pkt_r_instr__29_, issue_pkt_r_instr__28_, issue_pkt_r_instr__27_, issue_pkt_r_instr__26_, issue_pkt_r_instr__25_, issue_pkt_r_instr__24_, issue_pkt_r_instr__23_, issue_pkt_r_instr__22_, issue_pkt_r_instr__21_, issue_pkt_r_instr__20_, issue_pkt_r_instr__19_, issue_pkt_r_instr__18_, issue_pkt_r_instr__17_, issue_pkt_r_instr__16_, issue_pkt_r_instr__15_, issue_pkt_r_instr__14_, issue_pkt_r_instr__13_, issue_pkt_r_instr__12_, issue_pkt_r_instr__11_, issue_pkt_r_instr__10_, issue_pkt_r_instr__9_, issue_pkt_r_instr__8_, issue_pkt_r_instr__7_, issue_pkt_r_instr__6_, issue_pkt_r_instr__5_, issue_pkt_r_instr__4_, issue_pkt_r_instr__3_, issue_pkt_r_instr__2_, issue_pkt_r_instr__1_, issue_pkt_r_instr__0_, calc_status_o[236:236], calc_status_o[229:229], calc_status_o[235:235], calc_status_o[228:228], calc_status_o[234:230], calc_status_o[227:223], dispatch_pkt_instr_operands__imm__63_, dispatch_pkt_instr_operands__imm__62_, dispatch_pkt_instr_operands__imm__61_, dispatch_pkt_instr_operands__imm__60_, dispatch_pkt_instr_operands__imm__59_, dispatch_pkt_instr_operands__imm__58_, dispatch_pkt_instr_operands__imm__57_, dispatch_pkt_instr_operands__imm__56_, dispatch_pkt_instr_operands__imm__55_, dispatch_pkt_instr_operands__imm__54_, dispatch_pkt_instr_operands__imm__53_, dispatch_pkt_instr_operands__imm__52_, dispatch_pkt_instr_operands__imm__51_, dispatch_pkt_instr_operands__imm__50_, dispatch_pkt_instr_operands__imm__49_, dispatch_pkt_instr_operands__imm__48_, dispatch_pkt_instr_operands__imm__47_, dispatch_pkt_instr_operands__imm__46_, dispatch_pkt_instr_operands__imm__45_, dispatch_pkt_instr_operands__imm__44_, dispatch_pkt_instr_operands__imm__43_, dispatch_pkt_instr_operands__imm__42_, dispatch_pkt_instr_operands__imm__41_, dispatch_pkt_instr_operands__imm__40_, dispatch_pkt_instr_operands__imm__39_, dispatch_pkt_instr_operands__imm__38_, dispatch_pkt_instr_operands__imm__37_, dispatch_pkt_instr_operands__imm__36_, dispatch_pkt_instr_operands__imm__35_, dispatch_pkt_instr_operands__imm__34_, dispatch_pkt_instr_operands__imm__33_, dispatch_pkt_instr_operands__imm__32_, dispatch_pkt_instr_operands__imm__31_, dispatch_pkt_instr_operands__imm__30_, dispatch_pkt_instr_operands__imm__29_, dispatch_pkt_instr_operands__imm__28_, dispatch_pkt_instr_operands__imm__27_, dispatch_pkt_instr_operands__imm__26_, dispatch_pkt_instr_operands__imm__25_, dispatch_pkt_instr_operands__imm__24_, dispatch_pkt_instr_operands__imm__23_, dispatch_pkt_instr_operands__imm__22_, dispatch_pkt_instr_operands__imm__21_, dispatch_pkt_instr_operands__imm__20_, dispatch_pkt_instr_operands__imm__19_, dispatch_pkt_instr_operands__imm__18_, dispatch_pkt_instr_operands__imm__17_, dispatch_pkt_instr_operands__imm__16_, dispatch_pkt_instr_operands__imm__15_, dispatch_pkt_instr_operands__imm__14_, dispatch_pkt_instr_operands__imm__13_, dispatch_pkt_instr_operands__imm__12_, dispatch_pkt_instr_operands__imm__11_, dispatch_pkt_instr_operands__imm__10_, dispatch_pkt_instr_operands__imm__9_, dispatch_pkt_instr_operands__imm__8_, dispatch_pkt_instr_operands__imm__7_, dispatch_pkt_instr_operands__imm__6_, dispatch_pkt_instr_operands__imm__5_, dispatch_pkt_instr_operands__imm__4_, dispatch_pkt_instr_operands__imm__3_, dispatch_pkt_instr_operands__imm__2_, dispatch_pkt_instr_operands__imm__1_, dispatch_pkt_instr_operands__imm__0_ })
  );


  bsg_dff_reset_en_width_p1
  issue_v_reg
  (
    .clk_i(clk_i),
    .reset_i(n_16_net_),
    .en_i(n_17_net_),
    .data_i(issue_pkt_v_i),
    .data_o(calc_status_o[301])
  );


  bp_be_instr_decoder
  instr_decoder
  (
    .instr_i({ issue_pkt_r_instr__31_, issue_pkt_r_instr__30_, issue_pkt_r_instr__29_, issue_pkt_r_instr__28_, issue_pkt_r_instr__27_, issue_pkt_r_instr__26_, issue_pkt_r_instr__25_, issue_pkt_r_instr__24_, issue_pkt_r_instr__23_, issue_pkt_r_instr__22_, issue_pkt_r_instr__21_, issue_pkt_r_instr__20_, issue_pkt_r_instr__19_, issue_pkt_r_instr__18_, issue_pkt_r_instr__17_, issue_pkt_r_instr__16_, issue_pkt_r_instr__15_, issue_pkt_r_instr__14_, issue_pkt_r_instr__13_, issue_pkt_r_instr__12_, issue_pkt_r_instr__11_, issue_pkt_r_instr__10_, issue_pkt_r_instr__9_, issue_pkt_r_instr__8_, issue_pkt_r_instr__7_, issue_pkt_r_instr__6_, issue_pkt_r_instr__5_, issue_pkt_r_instr__4_, issue_pkt_r_instr__3_, issue_pkt_r_instr__2_, issue_pkt_r_instr__1_, issue_pkt_r_instr__0_ }),
    .fe_nop_v_i(n_18_net_),
    .be_nop_v_i(n_19_net_),
    .me_nop_v_i(n_20_net_),
    .decode_o({ dispatch_pkt_decode__instr_v_, dispatch_pkt_decode__fe_nop_v_, dispatch_pkt_decode__be_nop_v_, dispatch_pkt_decode__me_nop_v_, dispatch_pkt_decode__pipe_comp_v_, dispatch_pkt_decode__pipe_int_v_, dispatch_pkt_decode__pipe_mul_v_, dispatch_pkt_decode__pipe_mem_v_, dispatch_pkt_decode__pipe_fp_v_, dispatch_pkt_decode__irf_w_v_, dispatch_pkt_decode__frf_w_v_, dispatch_pkt_decode__mhartid_r_v_, dispatch_pkt_decode__dcache_w_v_, dispatch_pkt_decode__dcache_r_v_, decoded_fp_not_int_v_, dispatch_pkt_decode__ret_v_, dispatch_pkt_decode__amo_v_, dispatch_pkt_decode__jmp_v_, dispatch_pkt_decode__br_v_, dispatch_pkt_decode__opw_v_, decoded_fu_op_o, decoded_rs1_addr__4_, decoded_rs1_addr__3_, decoded_rs1_addr__2_, decoded_rs1_addr__1_, decoded_rs1_addr__0_, decoded_rs2_addr__4_, decoded_rs2_addr__3_, decoded_rs2_addr__2_, decoded_rs2_addr__1_, decoded_rs2_addr__0_, dispatch_pkt_decode__rd_addr__4_, dispatch_pkt_decode__rd_addr__3_, dispatch_pkt_decode__rd_addr__2_, dispatch_pkt_decode__rd_addr__1_, dispatch_pkt_decode__rd_addr__0_, dispatch_pkt_decode__src1_sel_, dispatch_pkt_decode__src2_sel_, dispatch_pkt_decode__baddr_sel_, dispatch_pkt_decode__result_sel_ }),
    .illegal_instr_o(exc_stage_n_0__illegal_instr_v_)
  );


  bp_be_bypass_fwd_els_p4
  int_bypass
  (
    .id_rs1_v_i(calc_status_o[236]),
    .id_rs1_addr_i({ decoded_rs1_addr__4_, decoded_rs1_addr__3_, decoded_rs1_addr__2_, decoded_rs1_addr__1_, decoded_rs1_addr__0_ }),
    .id_rs1_i(irf_rs1),
    .id_rs2_v_i(calc_status_o[229]),
    .id_rs2_addr_i({ decoded_rs2_addr__4_, decoded_rs2_addr__3_, decoded_rs2_addr__2_, decoded_rs2_addr__1_, decoded_rs2_addr__0_ }),
    .id_rs2_i(irf_rs2),
    .fwd_rd_v_i(comp_stage_n_slice_iwb_v),
    .fwd_rd_addr_i({ calc_status_o[103:99], calc_status_o[93:89], calc_status_o[83:79], calc_status_o[73:69] }),
    .fwd_rd_i({ comp_stage_n[639:576], comp_stage_n[511:448], comp_stage_n[383:320], comp_stage_n[255:192] }),
    .bypass_rs1_o(bypass_irs1),
    .bypass_rs2_o(bypass_irs2)
  );


  bp_be_bypass_fwd_els_p4
  fp_bypass
  (
    .id_rs1_v_i(calc_status_o[235]),
    .id_rs1_addr_i({ decoded_rs1_addr__4_, decoded_rs1_addr__3_, decoded_rs1_addr__2_, decoded_rs1_addr__1_, decoded_rs1_addr__0_ }),
    .id_rs1_i(frf_rs1),
    .id_rs2_v_i(calc_status_o[228]),
    .id_rs2_addr_i({ decoded_rs2_addr__4_, decoded_rs2_addr__3_, decoded_rs2_addr__2_, decoded_rs2_addr__1_, decoded_rs2_addr__0_ }),
    .id_rs2_i(frf_rs2),
    .fwd_rd_v_i(comp_stage_n_slice_fwb_v),
    .fwd_rd_addr_i({ calc_status_o[103:99], calc_status_o[93:89], calc_status_o[83:79], calc_status_o[73:69] }),
    .fwd_rd_i({ comp_stage_n[639:576], comp_stage_n[511:448], comp_stage_n[383:320], comp_stage_n[255:192] }),
    .bypass_rs1_o(bypass_frs1),
    .bypass_rs2_o(bypass_frs2)
  );


  bsg_mux_width_p64_els_p2
  bypass_xrs1_mux
  (
    .data_i({ bypass_frs1, bypass_irs1 }),
    .sel_i(decoded_fp_not_int_v_),
    .data_o({ dispatch_pkt_instr_operands__rs1__63_, dispatch_pkt_instr_operands__rs1__62_, dispatch_pkt_instr_operands__rs1__61_, dispatch_pkt_instr_operands__rs1__60_, dispatch_pkt_instr_operands__rs1__59_, dispatch_pkt_instr_operands__rs1__58_, dispatch_pkt_instr_operands__rs1__57_, dispatch_pkt_instr_operands__rs1__56_, dispatch_pkt_instr_operands__rs1__55_, dispatch_pkt_instr_operands__rs1__54_, dispatch_pkt_instr_operands__rs1__53_, dispatch_pkt_instr_operands__rs1__52_, dispatch_pkt_instr_operands__rs1__51_, dispatch_pkt_instr_operands__rs1__50_, dispatch_pkt_instr_operands__rs1__49_, dispatch_pkt_instr_operands__rs1__48_, dispatch_pkt_instr_operands__rs1__47_, dispatch_pkt_instr_operands__rs1__46_, dispatch_pkt_instr_operands__rs1__45_, dispatch_pkt_instr_operands__rs1__44_, dispatch_pkt_instr_operands__rs1__43_, dispatch_pkt_instr_operands__rs1__42_, dispatch_pkt_instr_operands__rs1__41_, dispatch_pkt_instr_operands__rs1__40_, dispatch_pkt_instr_operands__rs1__39_, dispatch_pkt_instr_operands__rs1__38_, dispatch_pkt_instr_operands__rs1__37_, dispatch_pkt_instr_operands__rs1__36_, dispatch_pkt_instr_operands__rs1__35_, dispatch_pkt_instr_operands__rs1__34_, dispatch_pkt_instr_operands__rs1__33_, dispatch_pkt_instr_operands__rs1__32_, dispatch_pkt_instr_operands__rs1__31_, dispatch_pkt_instr_operands__rs1__30_, dispatch_pkt_instr_operands__rs1__29_, dispatch_pkt_instr_operands__rs1__28_, dispatch_pkt_instr_operands__rs1__27_, dispatch_pkt_instr_operands__rs1__26_, dispatch_pkt_instr_operands__rs1__25_, dispatch_pkt_instr_operands__rs1__24_, dispatch_pkt_instr_operands__rs1__23_, dispatch_pkt_instr_operands__rs1__22_, dispatch_pkt_instr_operands__rs1__21_, dispatch_pkt_instr_operands__rs1__20_, dispatch_pkt_instr_operands__rs1__19_, dispatch_pkt_instr_operands__rs1__18_, dispatch_pkt_instr_operands__rs1__17_, dispatch_pkt_instr_operands__rs1__16_, dispatch_pkt_instr_operands__rs1__15_, dispatch_pkt_instr_operands__rs1__14_, dispatch_pkt_instr_operands__rs1__13_, dispatch_pkt_instr_operands__rs1__12_, dispatch_pkt_instr_operands__rs1__11_, dispatch_pkt_instr_operands__rs1__10_, dispatch_pkt_instr_operands__rs1__9_, dispatch_pkt_instr_operands__rs1__8_, dispatch_pkt_instr_operands__rs1__7_, dispatch_pkt_instr_operands__rs1__6_, dispatch_pkt_instr_operands__rs1__5_, dispatch_pkt_instr_operands__rs1__4_, dispatch_pkt_instr_operands__rs1__3_, dispatch_pkt_instr_operands__rs1__2_, dispatch_pkt_instr_operands__rs1__1_, dispatch_pkt_instr_operands__rs1__0_ })
  );


  bsg_mux_width_p64_els_p2
  bypass_xrs2_mux
  (
    .data_i({ bypass_frs2, bypass_irs2 }),
    .sel_i(decoded_fp_not_int_v_),
    .data_o({ dispatch_pkt_instr_operands__rs2__63_, dispatch_pkt_instr_operands__rs2__62_, dispatch_pkt_instr_operands__rs2__61_, dispatch_pkt_instr_operands__rs2__60_, dispatch_pkt_instr_operands__rs2__59_, dispatch_pkt_instr_operands__rs2__58_, dispatch_pkt_instr_operands__rs2__57_, dispatch_pkt_instr_operands__rs2__56_, dispatch_pkt_instr_operands__rs2__55_, dispatch_pkt_instr_operands__rs2__54_, dispatch_pkt_instr_operands__rs2__53_, dispatch_pkt_instr_operands__rs2__52_, dispatch_pkt_instr_operands__rs2__51_, dispatch_pkt_instr_operands__rs2__50_, dispatch_pkt_instr_operands__rs2__49_, dispatch_pkt_instr_operands__rs2__48_, dispatch_pkt_instr_operands__rs2__47_, dispatch_pkt_instr_operands__rs2__46_, dispatch_pkt_instr_operands__rs2__45_, dispatch_pkt_instr_operands__rs2__44_, dispatch_pkt_instr_operands__rs2__43_, dispatch_pkt_instr_operands__rs2__42_, dispatch_pkt_instr_operands__rs2__41_, dispatch_pkt_instr_operands__rs2__40_, dispatch_pkt_instr_operands__rs2__39_, dispatch_pkt_instr_operands__rs2__38_, dispatch_pkt_instr_operands__rs2__37_, dispatch_pkt_instr_operands__rs2__36_, dispatch_pkt_instr_operands__rs2__35_, dispatch_pkt_instr_operands__rs2__34_, dispatch_pkt_instr_operands__rs2__33_, dispatch_pkt_instr_operands__rs2__32_, dispatch_pkt_instr_operands__rs2__31_, dispatch_pkt_instr_operands__rs2__30_, dispatch_pkt_instr_operands__rs2__29_, dispatch_pkt_instr_operands__rs2__28_, dispatch_pkt_instr_operands__rs2__27_, dispatch_pkt_instr_operands__rs2__26_, dispatch_pkt_instr_operands__rs2__25_, dispatch_pkt_instr_operands__rs2__24_, dispatch_pkt_instr_operands__rs2__23_, dispatch_pkt_instr_operands__rs2__22_, dispatch_pkt_instr_operands__rs2__21_, dispatch_pkt_instr_operands__rs2__20_, dispatch_pkt_instr_operands__rs2__19_, dispatch_pkt_instr_operands__rs2__18_, dispatch_pkt_instr_operands__rs2__17_, dispatch_pkt_instr_operands__rs2__16_, dispatch_pkt_instr_operands__rs2__15_, dispatch_pkt_instr_operands__rs2__14_, dispatch_pkt_instr_operands__rs2__13_, dispatch_pkt_instr_operands__rs2__12_, dispatch_pkt_instr_operands__rs2__11_, dispatch_pkt_instr_operands__rs2__10_, dispatch_pkt_instr_operands__rs2__9_, dispatch_pkt_instr_operands__rs2__8_, dispatch_pkt_instr_operands__rs2__7_, dispatch_pkt_instr_operands__rs2__6_, dispatch_pkt_instr_operands__rs2__5_, dispatch_pkt_instr_operands__rs2__4_, dispatch_pkt_instr_operands__rs2__3_, dispatch_pkt_instr_operands__rs2__2_, dispatch_pkt_instr_operands__rs2__1_, dispatch_pkt_instr_operands__rs2__0_ })
  );


  bp_be_pipe_int_core_els_p1
  pipe_int
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .decode_i({ calc_stage_r_0__decode__instr_v_, calc_stage_r_0__decode__fe_nop_v_, calc_stage_r_0__decode__be_nop_v_, calc_stage_r_0__decode__me_nop_v_, calc_stage_r_0__decode__pipe_comp_v_, calc_stage_r_0__decode__pipe_int_v_, calc_stage_r_0__decode__pipe_mul_v_, calc_stage_r_0__decode__pipe_mem_v_, calc_stage_r_0__decode__pipe_fp_v_, calc_stage_r_0__decode__irf_w_v_, calc_stage_r_0__decode__frf_w_v_, calc_stage_r_0__decode__mhartid_r_v_, calc_stage_r_0__decode__dcache_w_v_, calc_stage_r_0__decode__dcache_r_v_, calc_stage_r_0__decode__fp_not_int_v_, calc_stage_r_0__decode__ret_v_, calc_stage_r_0__decode__amo_v_, calc_stage_r_0__decode__jmp_v_, calc_stage_r_0__decode__br_v_, calc_stage_r_0__decode__opw_v_, calc_stage_r_0__decode__fu_op__fu_op__3_, calc_stage_r_0__decode__fu_op__fu_op__2_, calc_stage_r_0__decode__fu_op__fu_op__1_, calc_stage_r_0__decode__fu_op__fu_op__0_, calc_stage_r_0__decode__rs1_addr__4_, calc_stage_r_0__decode__rs1_addr__3_, calc_stage_r_0__decode__rs1_addr__2_, calc_stage_r_0__decode__rs1_addr__1_, calc_stage_r_0__decode__rs1_addr__0_, calc_stage_r_0__decode__rs2_addr__4_, calc_stage_r_0__decode__rs2_addr__3_, calc_stage_r_0__decode__rs2_addr__2_, calc_stage_r_0__decode__rs2_addr__1_, calc_stage_r_0__decode__rs2_addr__0_, calc_status_o[73:69], calc_stage_r_0__decode__src1_sel_, calc_stage_r_0__decode__src2_sel_, calc_stage_r_0__decode__baddr_sel_, calc_stage_r_0__decode__result_sel_ }),
    .pc_i({ calc_stage_r_0__instr_metadata__pc__63_, calc_stage_r_0__instr_metadata__pc__62_, calc_stage_r_0__instr_metadata__pc__61_, calc_stage_r_0__instr_metadata__pc__60_, calc_stage_r_0__instr_metadata__pc__59_, calc_stage_r_0__instr_metadata__pc__58_, calc_stage_r_0__instr_metadata__pc__57_, calc_stage_r_0__instr_metadata__pc__56_, calc_stage_r_0__instr_metadata__pc__55_, calc_stage_r_0__instr_metadata__pc__54_, calc_stage_r_0__instr_metadata__pc__53_, calc_stage_r_0__instr_metadata__pc__52_, calc_stage_r_0__instr_metadata__pc__51_, calc_stage_r_0__instr_metadata__pc__50_, calc_stage_r_0__instr_metadata__pc__49_, calc_stage_r_0__instr_metadata__pc__48_, calc_stage_r_0__instr_metadata__pc__47_, calc_stage_r_0__instr_metadata__pc__46_, calc_stage_r_0__instr_metadata__pc__45_, calc_stage_r_0__instr_metadata__pc__44_, calc_stage_r_0__instr_metadata__pc__43_, calc_stage_r_0__instr_metadata__pc__42_, calc_stage_r_0__instr_metadata__pc__41_, calc_stage_r_0__instr_metadata__pc__40_, calc_stage_r_0__instr_metadata__pc__39_, calc_stage_r_0__instr_metadata__pc__38_, calc_stage_r_0__instr_metadata__pc__37_, calc_stage_r_0__instr_metadata__pc__36_, calc_stage_r_0__instr_metadata__pc__35_, calc_stage_r_0__instr_metadata__pc__34_, calc_stage_r_0__instr_metadata__pc__33_, calc_stage_r_0__instr_metadata__pc__32_, calc_stage_r_0__instr_metadata__pc__31_, calc_stage_r_0__instr_metadata__pc__30_, calc_stage_r_0__instr_metadata__pc__29_, calc_stage_r_0__instr_metadata__pc__28_, calc_stage_r_0__instr_metadata__pc__27_, calc_stage_r_0__instr_metadata__pc__26_, calc_stage_r_0__instr_metadata__pc__25_, calc_stage_r_0__instr_metadata__pc__24_, calc_stage_r_0__instr_metadata__pc__23_, calc_stage_r_0__instr_metadata__pc__22_, calc_stage_r_0__instr_metadata__pc__21_, calc_stage_r_0__instr_metadata__pc__20_, calc_stage_r_0__instr_metadata__pc__19_, calc_stage_r_0__instr_metadata__pc__18_, calc_stage_r_0__instr_metadata__pc__17_, calc_stage_r_0__instr_metadata__pc__16_, calc_stage_r_0__instr_metadata__pc__15_, calc_stage_r_0__instr_metadata__pc__14_, calc_stage_r_0__instr_metadata__pc__13_, calc_stage_r_0__instr_metadata__pc__12_, calc_stage_r_0__instr_metadata__pc__11_, calc_stage_r_0__instr_metadata__pc__10_, calc_stage_r_0__instr_metadata__pc__9_, calc_stage_r_0__instr_metadata__pc__8_, calc_stage_r_0__instr_metadata__pc__7_, calc_stage_r_0__instr_metadata__pc__6_, calc_stage_r_0__instr_metadata__pc__5_, calc_stage_r_0__instr_metadata__pc__4_, calc_stage_r_0__instr_metadata__pc__3_, calc_stage_r_0__instr_metadata__pc__2_, calc_stage_r_0__instr_metadata__pc__1_, calc_stage_r_0__instr_metadata__pc__0_ }),
    .rs1_i({ calc_stage_r_0__instr_operands__rs1__63_, calc_stage_r_0__instr_operands__rs1__62_, calc_stage_r_0__instr_operands__rs1__61_, calc_stage_r_0__instr_operands__rs1__60_, calc_stage_r_0__instr_operands__rs1__59_, calc_stage_r_0__instr_operands__rs1__58_, calc_stage_r_0__instr_operands__rs1__57_, calc_stage_r_0__instr_operands__rs1__56_, calc_stage_r_0__instr_operands__rs1__55_, calc_stage_r_0__instr_operands__rs1__54_, calc_stage_r_0__instr_operands__rs1__53_, calc_stage_r_0__instr_operands__rs1__52_, calc_stage_r_0__instr_operands__rs1__51_, calc_stage_r_0__instr_operands__rs1__50_, calc_stage_r_0__instr_operands__rs1__49_, calc_stage_r_0__instr_operands__rs1__48_, calc_stage_r_0__instr_operands__rs1__47_, calc_stage_r_0__instr_operands__rs1__46_, calc_stage_r_0__instr_operands__rs1__45_, calc_stage_r_0__instr_operands__rs1__44_, calc_stage_r_0__instr_operands__rs1__43_, calc_stage_r_0__instr_operands__rs1__42_, calc_stage_r_0__instr_operands__rs1__41_, calc_stage_r_0__instr_operands__rs1__40_, calc_stage_r_0__instr_operands__rs1__39_, calc_stage_r_0__instr_operands__rs1__38_, calc_stage_r_0__instr_operands__rs1__37_, calc_stage_r_0__instr_operands__rs1__36_, calc_stage_r_0__instr_operands__rs1__35_, calc_stage_r_0__instr_operands__rs1__34_, calc_stage_r_0__instr_operands__rs1__33_, calc_stage_r_0__instr_operands__rs1__32_, calc_stage_r_0__instr_operands__rs1__31_, calc_stage_r_0__instr_operands__rs1__30_, calc_stage_r_0__instr_operands__rs1__29_, calc_stage_r_0__instr_operands__rs1__28_, calc_stage_r_0__instr_operands__rs1__27_, calc_stage_r_0__instr_operands__rs1__26_, calc_stage_r_0__instr_operands__rs1__25_, calc_stage_r_0__instr_operands__rs1__24_, calc_stage_r_0__instr_operands__rs1__23_, calc_stage_r_0__instr_operands__rs1__22_, calc_stage_r_0__instr_operands__rs1__21_, calc_stage_r_0__instr_operands__rs1__20_, calc_stage_r_0__instr_operands__rs1__19_, calc_stage_r_0__instr_operands__rs1__18_, calc_stage_r_0__instr_operands__rs1__17_, calc_stage_r_0__instr_operands__rs1__16_, calc_stage_r_0__instr_operands__rs1__15_, calc_stage_r_0__instr_operands__rs1__14_, calc_stage_r_0__instr_operands__rs1__13_, calc_stage_r_0__instr_operands__rs1__12_, calc_stage_r_0__instr_operands__rs1__11_, calc_stage_r_0__instr_operands__rs1__10_, calc_stage_r_0__instr_operands__rs1__9_, calc_stage_r_0__instr_operands__rs1__8_, calc_stage_r_0__instr_operands__rs1__7_, calc_stage_r_0__instr_operands__rs1__6_, calc_stage_r_0__instr_operands__rs1__5_, calc_stage_r_0__instr_operands__rs1__4_, calc_stage_r_0__instr_operands__rs1__3_, calc_stage_r_0__instr_operands__rs1__2_, calc_stage_r_0__instr_operands__rs1__1_, calc_stage_r_0__instr_operands__rs1__0_ }),
    .rs2_i({ calc_stage_r_0__instr_operands__rs2__63_, calc_stage_r_0__instr_operands__rs2__62_, calc_stage_r_0__instr_operands__rs2__61_, calc_stage_r_0__instr_operands__rs2__60_, calc_stage_r_0__instr_operands__rs2__59_, calc_stage_r_0__instr_operands__rs2__58_, calc_stage_r_0__instr_operands__rs2__57_, calc_stage_r_0__instr_operands__rs2__56_, calc_stage_r_0__instr_operands__rs2__55_, calc_stage_r_0__instr_operands__rs2__54_, calc_stage_r_0__instr_operands__rs2__53_, calc_stage_r_0__instr_operands__rs2__52_, calc_stage_r_0__instr_operands__rs2__51_, calc_stage_r_0__instr_operands__rs2__50_, calc_stage_r_0__instr_operands__rs2__49_, calc_stage_r_0__instr_operands__rs2__48_, calc_stage_r_0__instr_operands__rs2__47_, calc_stage_r_0__instr_operands__rs2__46_, calc_stage_r_0__instr_operands__rs2__45_, calc_stage_r_0__instr_operands__rs2__44_, calc_stage_r_0__instr_operands__rs2__43_, calc_stage_r_0__instr_operands__rs2__42_, calc_stage_r_0__instr_operands__rs2__41_, calc_stage_r_0__instr_operands__rs2__40_, calc_stage_r_0__instr_operands__rs2__39_, calc_stage_r_0__instr_operands__rs2__38_, calc_stage_r_0__instr_operands__rs2__37_, calc_stage_r_0__instr_operands__rs2__36_, calc_stage_r_0__instr_operands__rs2__35_, calc_stage_r_0__instr_operands__rs2__34_, calc_stage_r_0__instr_operands__rs2__33_, calc_stage_r_0__instr_operands__rs2__32_, calc_stage_r_0__instr_operands__rs2__31_, calc_stage_r_0__instr_operands__rs2__30_, calc_stage_r_0__instr_operands__rs2__29_, calc_stage_r_0__instr_operands__rs2__28_, calc_stage_r_0__instr_operands__rs2__27_, calc_stage_r_0__instr_operands__rs2__26_, calc_stage_r_0__instr_operands__rs2__25_, calc_stage_r_0__instr_operands__rs2__24_, calc_stage_r_0__instr_operands__rs2__23_, calc_stage_r_0__instr_operands__rs2__22_, calc_stage_r_0__instr_operands__rs2__21_, calc_stage_r_0__instr_operands__rs2__20_, calc_stage_r_0__instr_operands__rs2__19_, calc_stage_r_0__instr_operands__rs2__18_, calc_stage_r_0__instr_operands__rs2__17_, calc_stage_r_0__instr_operands__rs2__16_, calc_stage_r_0__instr_operands__rs2__15_, calc_stage_r_0__instr_operands__rs2__14_, calc_stage_r_0__instr_operands__rs2__13_, calc_stage_r_0__instr_operands__rs2__12_, calc_stage_r_0__instr_operands__rs2__11_, calc_stage_r_0__instr_operands__rs2__10_, calc_stage_r_0__instr_operands__rs2__9_, calc_stage_r_0__instr_operands__rs2__8_, calc_stage_r_0__instr_operands__rs2__7_, calc_stage_r_0__instr_operands__rs2__6_, calc_stage_r_0__instr_operands__rs2__5_, calc_stage_r_0__instr_operands__rs2__4_, calc_stage_r_0__instr_operands__rs2__3_, calc_stage_r_0__instr_operands__rs2__2_, calc_stage_r_0__instr_operands__rs2__1_, calc_stage_r_0__instr_operands__rs2__0_ }),
    .imm_i({ calc_stage_r_0__instr_operands__imm__63_, calc_stage_r_0__instr_operands__imm__62_, calc_stage_r_0__instr_operands__imm__61_, calc_stage_r_0__instr_operands__imm__60_, calc_stage_r_0__instr_operands__imm__59_, calc_stage_r_0__instr_operands__imm__58_, calc_stage_r_0__instr_operands__imm__57_, calc_stage_r_0__instr_operands__imm__56_, calc_stage_r_0__instr_operands__imm__55_, calc_stage_r_0__instr_operands__imm__54_, calc_stage_r_0__instr_operands__imm__53_, calc_stage_r_0__instr_operands__imm__52_, calc_stage_r_0__instr_operands__imm__51_, calc_stage_r_0__instr_operands__imm__50_, calc_stage_r_0__instr_operands__imm__49_, calc_stage_r_0__instr_operands__imm__48_, calc_stage_r_0__instr_operands__imm__47_, calc_stage_r_0__instr_operands__imm__46_, calc_stage_r_0__instr_operands__imm__45_, calc_stage_r_0__instr_operands__imm__44_, calc_stage_r_0__instr_operands__imm__43_, calc_stage_r_0__instr_operands__imm__42_, calc_stage_r_0__instr_operands__imm__41_, calc_stage_r_0__instr_operands__imm__40_, calc_stage_r_0__instr_operands__imm__39_, calc_stage_r_0__instr_operands__imm__38_, calc_stage_r_0__instr_operands__imm__37_, calc_stage_r_0__instr_operands__imm__36_, calc_stage_r_0__instr_operands__imm__35_, calc_stage_r_0__instr_operands__imm__34_, calc_stage_r_0__instr_operands__imm__33_, calc_stage_r_0__instr_operands__imm__32_, calc_stage_r_0__instr_operands__imm__31_, calc_stage_r_0__instr_operands__imm__30_, calc_stage_r_0__instr_operands__imm__29_, calc_stage_r_0__instr_operands__imm__28_, calc_stage_r_0__instr_operands__imm__27_, calc_stage_r_0__instr_operands__imm__26_, calc_stage_r_0__instr_operands__imm__25_, calc_stage_r_0__instr_operands__imm__24_, calc_stage_r_0__instr_operands__imm__23_, calc_stage_r_0__instr_operands__imm__22_, calc_stage_r_0__instr_operands__imm__21_, calc_stage_r_0__instr_operands__imm__20_, calc_stage_r_0__instr_operands__imm__19_, calc_stage_r_0__instr_operands__imm__18_, calc_stage_r_0__instr_operands__imm__17_, calc_stage_r_0__instr_operands__imm__16_, calc_stage_r_0__instr_operands__imm__15_, calc_stage_r_0__instr_operands__imm__14_, calc_stage_r_0__instr_operands__imm__13_, calc_stage_r_0__instr_operands__imm__12_, calc_stage_r_0__instr_operands__imm__11_, calc_stage_r_0__instr_operands__imm__10_, calc_stage_r_0__instr_operands__imm__9_, calc_stage_r_0__instr_operands__imm__8_, calc_stage_r_0__instr_operands__imm__7_, calc_stage_r_0__instr_operands__imm__6_, calc_stage_r_0__instr_operands__imm__5_, calc_stage_r_0__instr_operands__imm__4_, calc_stage_r_0__instr_operands__imm__3_, calc_stage_r_0__instr_operands__imm__2_, calc_stage_r_0__instr_operands__imm__1_, calc_stage_r_0__instr_operands__imm__0_ }),
    .exc_i({ exc_stage_r_0__poison_v_, exc_stage_r_0__roll_v_, exc_stage_r_0__illegal_instr_v_, exc_stage_r_0__tlb_miss_v_, exc_stage_r_0__load_fault_v_, exc_stage_r_0__store_fault_v_, exc_stage_r_0__cache_miss_v_ }),
    .mhartid_i(proc_cfg_i[2]),
    .result_o({ int_calc_result_result__63_, int_calc_result_result__62_, int_calc_result_result__61_, int_calc_result_result__60_, int_calc_result_result__59_, int_calc_result_result__58_, int_calc_result_result__57_, int_calc_result_result__56_, int_calc_result_result__55_, int_calc_result_result__54_, int_calc_result_result__53_, int_calc_result_result__52_, int_calc_result_result__51_, int_calc_result_result__50_, int_calc_result_result__49_, int_calc_result_result__48_, int_calc_result_result__47_, int_calc_result_result__46_, int_calc_result_result__45_, int_calc_result_result__44_, int_calc_result_result__43_, int_calc_result_result__42_, int_calc_result_result__41_, int_calc_result_result__40_, int_calc_result_result__39_, int_calc_result_result__38_, int_calc_result_result__37_, int_calc_result_result__36_, int_calc_result_result__35_, int_calc_result_result__34_, int_calc_result_result__33_, int_calc_result_result__32_, int_calc_result_result__31_, int_calc_result_result__30_, int_calc_result_result__29_, int_calc_result_result__28_, int_calc_result_result__27_, int_calc_result_result__26_, int_calc_result_result__25_, int_calc_result_result__24_, int_calc_result_result__23_, int_calc_result_result__22_, int_calc_result_result__21_, int_calc_result_result__20_, int_calc_result_result__19_, int_calc_result_result__18_, int_calc_result_result__17_, int_calc_result_result__16_, int_calc_result_result__15_, int_calc_result_result__14_, int_calc_result_result__13_, int_calc_result_result__12_, int_calc_result_result__11_, int_calc_result_result__10_, int_calc_result_result__9_, int_calc_result_result__8_, int_calc_result_result__7_, int_calc_result_result__6_, int_calc_result_result__5_, int_calc_result_result__4_, int_calc_result_result__3_, int_calc_result_result__2_, int_calc_result_result__1_, int_calc_result_result__0_ }),
    .br_tgt_o(calc_status_o[221:158])
  );


  bp_be_pipe_mul
  pipe_mul
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .decode_i({ calc_stage_r_0__decode__instr_v_, calc_stage_r_0__decode__fe_nop_v_, calc_stage_r_0__decode__be_nop_v_, calc_stage_r_0__decode__me_nop_v_, calc_stage_r_0__decode__pipe_comp_v_, calc_stage_r_0__decode__pipe_int_v_, calc_stage_r_0__decode__pipe_mul_v_, calc_stage_r_0__decode__pipe_mem_v_, calc_stage_r_0__decode__pipe_fp_v_, calc_stage_r_0__decode__irf_w_v_, calc_stage_r_0__decode__frf_w_v_, calc_stage_r_0__decode__mhartid_r_v_, calc_stage_r_0__decode__dcache_w_v_, calc_stage_r_0__decode__dcache_r_v_, calc_stage_r_0__decode__fp_not_int_v_, calc_stage_r_0__decode__ret_v_, calc_stage_r_0__decode__amo_v_, calc_stage_r_0__decode__jmp_v_, calc_stage_r_0__decode__br_v_, calc_stage_r_0__decode__opw_v_, calc_stage_r_0__decode__fu_op__fu_op__3_, calc_stage_r_0__decode__fu_op__fu_op__2_, calc_stage_r_0__decode__fu_op__fu_op__1_, calc_stage_r_0__decode__fu_op__fu_op__0_, calc_stage_r_0__decode__rs1_addr__4_, calc_stage_r_0__decode__rs1_addr__3_, calc_stage_r_0__decode__rs1_addr__2_, calc_stage_r_0__decode__rs1_addr__1_, calc_stage_r_0__decode__rs1_addr__0_, calc_stage_r_0__decode__rs2_addr__4_, calc_stage_r_0__decode__rs2_addr__3_, calc_stage_r_0__decode__rs2_addr__2_, calc_stage_r_0__decode__rs2_addr__1_, calc_stage_r_0__decode__rs2_addr__0_, calc_status_o[73:69], calc_stage_r_0__decode__src1_sel_, calc_stage_r_0__decode__src2_sel_, calc_stage_r_0__decode__baddr_sel_, calc_stage_r_0__decode__result_sel_ }),
    .rs1_i({ calc_stage_r_0__instr_operands__rs1__63_, calc_stage_r_0__instr_operands__rs1__62_, calc_stage_r_0__instr_operands__rs1__61_, calc_stage_r_0__instr_operands__rs1__60_, calc_stage_r_0__instr_operands__rs1__59_, calc_stage_r_0__instr_operands__rs1__58_, calc_stage_r_0__instr_operands__rs1__57_, calc_stage_r_0__instr_operands__rs1__56_, calc_stage_r_0__instr_operands__rs1__55_, calc_stage_r_0__instr_operands__rs1__54_, calc_stage_r_0__instr_operands__rs1__53_, calc_stage_r_0__instr_operands__rs1__52_, calc_stage_r_0__instr_operands__rs1__51_, calc_stage_r_0__instr_operands__rs1__50_, calc_stage_r_0__instr_operands__rs1__49_, calc_stage_r_0__instr_operands__rs1__48_, calc_stage_r_0__instr_operands__rs1__47_, calc_stage_r_0__instr_operands__rs1__46_, calc_stage_r_0__instr_operands__rs1__45_, calc_stage_r_0__instr_operands__rs1__44_, calc_stage_r_0__instr_operands__rs1__43_, calc_stage_r_0__instr_operands__rs1__42_, calc_stage_r_0__instr_operands__rs1__41_, calc_stage_r_0__instr_operands__rs1__40_, calc_stage_r_0__instr_operands__rs1__39_, calc_stage_r_0__instr_operands__rs1__38_, calc_stage_r_0__instr_operands__rs1__37_, calc_stage_r_0__instr_operands__rs1__36_, calc_stage_r_0__instr_operands__rs1__35_, calc_stage_r_0__instr_operands__rs1__34_, calc_stage_r_0__instr_operands__rs1__33_, calc_stage_r_0__instr_operands__rs1__32_, calc_stage_r_0__instr_operands__rs1__31_, calc_stage_r_0__instr_operands__rs1__30_, calc_stage_r_0__instr_operands__rs1__29_, calc_stage_r_0__instr_operands__rs1__28_, calc_stage_r_0__instr_operands__rs1__27_, calc_stage_r_0__instr_operands__rs1__26_, calc_stage_r_0__instr_operands__rs1__25_, calc_stage_r_0__instr_operands__rs1__24_, calc_stage_r_0__instr_operands__rs1__23_, calc_stage_r_0__instr_operands__rs1__22_, calc_stage_r_0__instr_operands__rs1__21_, calc_stage_r_0__instr_operands__rs1__20_, calc_stage_r_0__instr_operands__rs1__19_, calc_stage_r_0__instr_operands__rs1__18_, calc_stage_r_0__instr_operands__rs1__17_, calc_stage_r_0__instr_operands__rs1__16_, calc_stage_r_0__instr_operands__rs1__15_, calc_stage_r_0__instr_operands__rs1__14_, calc_stage_r_0__instr_operands__rs1__13_, calc_stage_r_0__instr_operands__rs1__12_, calc_stage_r_0__instr_operands__rs1__11_, calc_stage_r_0__instr_operands__rs1__10_, calc_stage_r_0__instr_operands__rs1__9_, calc_stage_r_0__instr_operands__rs1__8_, calc_stage_r_0__instr_operands__rs1__7_, calc_stage_r_0__instr_operands__rs1__6_, calc_stage_r_0__instr_operands__rs1__5_, calc_stage_r_0__instr_operands__rs1__4_, calc_stage_r_0__instr_operands__rs1__3_, calc_stage_r_0__instr_operands__rs1__2_, calc_stage_r_0__instr_operands__rs1__1_, calc_stage_r_0__instr_operands__rs1__0_ }),
    .rs2_i({ calc_stage_r_0__instr_operands__rs2__63_, calc_stage_r_0__instr_operands__rs2__62_, calc_stage_r_0__instr_operands__rs2__61_, calc_stage_r_0__instr_operands__rs2__60_, calc_stage_r_0__instr_operands__rs2__59_, calc_stage_r_0__instr_operands__rs2__58_, calc_stage_r_0__instr_operands__rs2__57_, calc_stage_r_0__instr_operands__rs2__56_, calc_stage_r_0__instr_operands__rs2__55_, calc_stage_r_0__instr_operands__rs2__54_, calc_stage_r_0__instr_operands__rs2__53_, calc_stage_r_0__instr_operands__rs2__52_, calc_stage_r_0__instr_operands__rs2__51_, calc_stage_r_0__instr_operands__rs2__50_, calc_stage_r_0__instr_operands__rs2__49_, calc_stage_r_0__instr_operands__rs2__48_, calc_stage_r_0__instr_operands__rs2__47_, calc_stage_r_0__instr_operands__rs2__46_, calc_stage_r_0__instr_operands__rs2__45_, calc_stage_r_0__instr_operands__rs2__44_, calc_stage_r_0__instr_operands__rs2__43_, calc_stage_r_0__instr_operands__rs2__42_, calc_stage_r_0__instr_operands__rs2__41_, calc_stage_r_0__instr_operands__rs2__40_, calc_stage_r_0__instr_operands__rs2__39_, calc_stage_r_0__instr_operands__rs2__38_, calc_stage_r_0__instr_operands__rs2__37_, calc_stage_r_0__instr_operands__rs2__36_, calc_stage_r_0__instr_operands__rs2__35_, calc_stage_r_0__instr_operands__rs2__34_, calc_stage_r_0__instr_operands__rs2__33_, calc_stage_r_0__instr_operands__rs2__32_, calc_stage_r_0__instr_operands__rs2__31_, calc_stage_r_0__instr_operands__rs2__30_, calc_stage_r_0__instr_operands__rs2__29_, calc_stage_r_0__instr_operands__rs2__28_, calc_stage_r_0__instr_operands__rs2__27_, calc_stage_r_0__instr_operands__rs2__26_, calc_stage_r_0__instr_operands__rs2__25_, calc_stage_r_0__instr_operands__rs2__24_, calc_stage_r_0__instr_operands__rs2__23_, calc_stage_r_0__instr_operands__rs2__22_, calc_stage_r_0__instr_operands__rs2__21_, calc_stage_r_0__instr_operands__rs2__20_, calc_stage_r_0__instr_operands__rs2__19_, calc_stage_r_0__instr_operands__rs2__18_, calc_stage_r_0__instr_operands__rs2__17_, calc_stage_r_0__instr_operands__rs2__16_, calc_stage_r_0__instr_operands__rs2__15_, calc_stage_r_0__instr_operands__rs2__14_, calc_stage_r_0__instr_operands__rs2__13_, calc_stage_r_0__instr_operands__rs2__12_, calc_stage_r_0__instr_operands__rs2__11_, calc_stage_r_0__instr_operands__rs2__10_, calc_stage_r_0__instr_operands__rs2__9_, calc_stage_r_0__instr_operands__rs2__8_, calc_stage_r_0__instr_operands__rs2__7_, calc_stage_r_0__instr_operands__rs2__6_, calc_stage_r_0__instr_operands__rs2__5_, calc_stage_r_0__instr_operands__rs2__4_, calc_stage_r_0__instr_operands__rs2__3_, calc_stage_r_0__instr_operands__rs2__2_, calc_stage_r_0__instr_operands__rs2__1_, calc_stage_r_0__instr_operands__rs2__0_ }),
    .exc_i({ exc_stage_r_0__poison_v_, exc_stage_r_0__roll_v_, exc_stage_r_0__illegal_instr_v_, exc_stage_r_0__tlb_miss_v_, exc_stage_r_0__load_fault_v_, exc_stage_r_0__store_fault_v_, exc_stage_r_0__cache_miss_v_ }),
    .result_o(mul_calc_result[127:64])
  );


  bp_be_pipe_mem_vaddr_width_p56_lce_sets_p64_cce_block_size_in_bytes_p64
  pipe_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .decode_i({ calc_stage_r_0__decode__instr_v_, calc_stage_r_0__decode__fe_nop_v_, calc_stage_r_0__decode__be_nop_v_, calc_stage_r_0__decode__me_nop_v_, calc_stage_r_0__decode__pipe_comp_v_, calc_stage_r_0__decode__pipe_int_v_, calc_stage_r_0__decode__pipe_mul_v_, calc_stage_r_0__decode__pipe_mem_v_, calc_stage_r_0__decode__pipe_fp_v_, calc_stage_r_0__decode__irf_w_v_, calc_stage_r_0__decode__frf_w_v_, calc_stage_r_0__decode__mhartid_r_v_, calc_stage_r_0__decode__dcache_w_v_, calc_stage_r_0__decode__dcache_r_v_, calc_stage_r_0__decode__fp_not_int_v_, calc_stage_r_0__decode__ret_v_, calc_stage_r_0__decode__amo_v_, calc_stage_r_0__decode__jmp_v_, calc_stage_r_0__decode__br_v_, calc_stage_r_0__decode__opw_v_, calc_stage_r_0__decode__fu_op__fu_op__3_, calc_stage_r_0__decode__fu_op__fu_op__2_, calc_stage_r_0__decode__fu_op__fu_op__1_, calc_stage_r_0__decode__fu_op__fu_op__0_, calc_stage_r_0__decode__rs1_addr__4_, calc_stage_r_0__decode__rs1_addr__3_, calc_stage_r_0__decode__rs1_addr__2_, calc_stage_r_0__decode__rs1_addr__1_, calc_stage_r_0__decode__rs1_addr__0_, calc_stage_r_0__decode__rs2_addr__4_, calc_stage_r_0__decode__rs2_addr__3_, calc_stage_r_0__decode__rs2_addr__2_, calc_stage_r_0__decode__rs2_addr__1_, calc_stage_r_0__decode__rs2_addr__0_, calc_status_o[73:69], calc_stage_r_0__decode__src1_sel_, calc_stage_r_0__decode__src2_sel_, calc_stage_r_0__decode__baddr_sel_, calc_stage_r_0__decode__result_sel_ }),
    .rs1_i({ calc_stage_r_0__instr_operands__rs1__63_, calc_stage_r_0__instr_operands__rs1__62_, calc_stage_r_0__instr_operands__rs1__61_, calc_stage_r_0__instr_operands__rs1__60_, calc_stage_r_0__instr_operands__rs1__59_, calc_stage_r_0__instr_operands__rs1__58_, calc_stage_r_0__instr_operands__rs1__57_, calc_stage_r_0__instr_operands__rs1__56_, calc_stage_r_0__instr_operands__rs1__55_, calc_stage_r_0__instr_operands__rs1__54_, calc_stage_r_0__instr_operands__rs1__53_, calc_stage_r_0__instr_operands__rs1__52_, calc_stage_r_0__instr_operands__rs1__51_, calc_stage_r_0__instr_operands__rs1__50_, calc_stage_r_0__instr_operands__rs1__49_, calc_stage_r_0__instr_operands__rs1__48_, calc_stage_r_0__instr_operands__rs1__47_, calc_stage_r_0__instr_operands__rs1__46_, calc_stage_r_0__instr_operands__rs1__45_, calc_stage_r_0__instr_operands__rs1__44_, calc_stage_r_0__instr_operands__rs1__43_, calc_stage_r_0__instr_operands__rs1__42_, calc_stage_r_0__instr_operands__rs1__41_, calc_stage_r_0__instr_operands__rs1__40_, calc_stage_r_0__instr_operands__rs1__39_, calc_stage_r_0__instr_operands__rs1__38_, calc_stage_r_0__instr_operands__rs1__37_, calc_stage_r_0__instr_operands__rs1__36_, calc_stage_r_0__instr_operands__rs1__35_, calc_stage_r_0__instr_operands__rs1__34_, calc_stage_r_0__instr_operands__rs1__33_, calc_stage_r_0__instr_operands__rs1__32_, calc_stage_r_0__instr_operands__rs1__31_, calc_stage_r_0__instr_operands__rs1__30_, calc_stage_r_0__instr_operands__rs1__29_, calc_stage_r_0__instr_operands__rs1__28_, calc_stage_r_0__instr_operands__rs1__27_, calc_stage_r_0__instr_operands__rs1__26_, calc_stage_r_0__instr_operands__rs1__25_, calc_stage_r_0__instr_operands__rs1__24_, calc_stage_r_0__instr_operands__rs1__23_, calc_stage_r_0__instr_operands__rs1__22_, calc_stage_r_0__instr_operands__rs1__21_, calc_stage_r_0__instr_operands__rs1__20_, calc_stage_r_0__instr_operands__rs1__19_, calc_stage_r_0__instr_operands__rs1__18_, calc_stage_r_0__instr_operands__rs1__17_, calc_stage_r_0__instr_operands__rs1__16_, calc_stage_r_0__instr_operands__rs1__15_, calc_stage_r_0__instr_operands__rs1__14_, calc_stage_r_0__instr_operands__rs1__13_, calc_stage_r_0__instr_operands__rs1__12_, calc_stage_r_0__instr_operands__rs1__11_, calc_stage_r_0__instr_operands__rs1__10_, calc_stage_r_0__instr_operands__rs1__9_, calc_stage_r_0__instr_operands__rs1__8_, calc_stage_r_0__instr_operands__rs1__7_, calc_stage_r_0__instr_operands__rs1__6_, calc_stage_r_0__instr_operands__rs1__5_, calc_stage_r_0__instr_operands__rs1__4_, calc_stage_r_0__instr_operands__rs1__3_, calc_stage_r_0__instr_operands__rs1__2_, calc_stage_r_0__instr_operands__rs1__1_, calc_stage_r_0__instr_operands__rs1__0_ }),
    .rs2_i({ calc_stage_r_0__instr_operands__rs2__63_, calc_stage_r_0__instr_operands__rs2__62_, calc_stage_r_0__instr_operands__rs2__61_, calc_stage_r_0__instr_operands__rs2__60_, calc_stage_r_0__instr_operands__rs2__59_, calc_stage_r_0__instr_operands__rs2__58_, calc_stage_r_0__instr_operands__rs2__57_, calc_stage_r_0__instr_operands__rs2__56_, calc_stage_r_0__instr_operands__rs2__55_, calc_stage_r_0__instr_operands__rs2__54_, calc_stage_r_0__instr_operands__rs2__53_, calc_stage_r_0__instr_operands__rs2__52_, calc_stage_r_0__instr_operands__rs2__51_, calc_stage_r_0__instr_operands__rs2__50_, calc_stage_r_0__instr_operands__rs2__49_, calc_stage_r_0__instr_operands__rs2__48_, calc_stage_r_0__instr_operands__rs2__47_, calc_stage_r_0__instr_operands__rs2__46_, calc_stage_r_0__instr_operands__rs2__45_, calc_stage_r_0__instr_operands__rs2__44_, calc_stage_r_0__instr_operands__rs2__43_, calc_stage_r_0__instr_operands__rs2__42_, calc_stage_r_0__instr_operands__rs2__41_, calc_stage_r_0__instr_operands__rs2__40_, calc_stage_r_0__instr_operands__rs2__39_, calc_stage_r_0__instr_operands__rs2__38_, calc_stage_r_0__instr_operands__rs2__37_, calc_stage_r_0__instr_operands__rs2__36_, calc_stage_r_0__instr_operands__rs2__35_, calc_stage_r_0__instr_operands__rs2__34_, calc_stage_r_0__instr_operands__rs2__33_, calc_stage_r_0__instr_operands__rs2__32_, calc_stage_r_0__instr_operands__rs2__31_, calc_stage_r_0__instr_operands__rs2__30_, calc_stage_r_0__instr_operands__rs2__29_, calc_stage_r_0__instr_operands__rs2__28_, calc_stage_r_0__instr_operands__rs2__27_, calc_stage_r_0__instr_operands__rs2__26_, calc_stage_r_0__instr_operands__rs2__25_, calc_stage_r_0__instr_operands__rs2__24_, calc_stage_r_0__instr_operands__rs2__23_, calc_stage_r_0__instr_operands__rs2__22_, calc_stage_r_0__instr_operands__rs2__21_, calc_stage_r_0__instr_operands__rs2__20_, calc_stage_r_0__instr_operands__rs2__19_, calc_stage_r_0__instr_operands__rs2__18_, calc_stage_r_0__instr_operands__rs2__17_, calc_stage_r_0__instr_operands__rs2__16_, calc_stage_r_0__instr_operands__rs2__15_, calc_stage_r_0__instr_operands__rs2__14_, calc_stage_r_0__instr_operands__rs2__13_, calc_stage_r_0__instr_operands__rs2__12_, calc_stage_r_0__instr_operands__rs2__11_, calc_stage_r_0__instr_operands__rs2__10_, calc_stage_r_0__instr_operands__rs2__9_, calc_stage_r_0__instr_operands__rs2__8_, calc_stage_r_0__instr_operands__rs2__7_, calc_stage_r_0__instr_operands__rs2__6_, calc_stage_r_0__instr_operands__rs2__5_, calc_stage_r_0__instr_operands__rs2__4_, calc_stage_r_0__instr_operands__rs2__3_, calc_stage_r_0__instr_operands__rs2__2_, calc_stage_r_0__instr_operands__rs2__1_, calc_stage_r_0__instr_operands__rs2__0_ }),
    .imm_i({ calc_stage_r_0__instr_operands__imm__63_, calc_stage_r_0__instr_operands__imm__62_, calc_stage_r_0__instr_operands__imm__61_, calc_stage_r_0__instr_operands__imm__60_, calc_stage_r_0__instr_operands__imm__59_, calc_stage_r_0__instr_operands__imm__58_, calc_stage_r_0__instr_operands__imm__57_, calc_stage_r_0__instr_operands__imm__56_, calc_stage_r_0__instr_operands__imm__55_, calc_stage_r_0__instr_operands__imm__54_, calc_stage_r_0__instr_operands__imm__53_, calc_stage_r_0__instr_operands__imm__52_, calc_stage_r_0__instr_operands__imm__51_, calc_stage_r_0__instr_operands__imm__50_, calc_stage_r_0__instr_operands__imm__49_, calc_stage_r_0__instr_operands__imm__48_, calc_stage_r_0__instr_operands__imm__47_, calc_stage_r_0__instr_operands__imm__46_, calc_stage_r_0__instr_operands__imm__45_, calc_stage_r_0__instr_operands__imm__44_, calc_stage_r_0__instr_operands__imm__43_, calc_stage_r_0__instr_operands__imm__42_, calc_stage_r_0__instr_operands__imm__41_, calc_stage_r_0__instr_operands__imm__40_, calc_stage_r_0__instr_operands__imm__39_, calc_stage_r_0__instr_operands__imm__38_, calc_stage_r_0__instr_operands__imm__37_, calc_stage_r_0__instr_operands__imm__36_, calc_stage_r_0__instr_operands__imm__35_, calc_stage_r_0__instr_operands__imm__34_, calc_stage_r_0__instr_operands__imm__33_, calc_stage_r_0__instr_operands__imm__32_, calc_stage_r_0__instr_operands__imm__31_, calc_stage_r_0__instr_operands__imm__30_, calc_stage_r_0__instr_operands__imm__29_, calc_stage_r_0__instr_operands__imm__28_, calc_stage_r_0__instr_operands__imm__27_, calc_stage_r_0__instr_operands__imm__26_, calc_stage_r_0__instr_operands__imm__25_, calc_stage_r_0__instr_operands__imm__24_, calc_stage_r_0__instr_operands__imm__23_, calc_stage_r_0__instr_operands__imm__22_, calc_stage_r_0__instr_operands__imm__21_, calc_stage_r_0__instr_operands__imm__20_, calc_stage_r_0__instr_operands__imm__19_, calc_stage_r_0__instr_operands__imm__18_, calc_stage_r_0__instr_operands__imm__17_, calc_stage_r_0__instr_operands__imm__16_, calc_stage_r_0__instr_operands__imm__15_, calc_stage_r_0__instr_operands__imm__14_, calc_stage_r_0__instr_operands__imm__13_, calc_stage_r_0__instr_operands__imm__12_, calc_stage_r_0__instr_operands__imm__11_, calc_stage_r_0__instr_operands__imm__10_, calc_stage_r_0__instr_operands__imm__9_, calc_stage_r_0__instr_operands__imm__8_, calc_stage_r_0__instr_operands__imm__7_, calc_stage_r_0__instr_operands__imm__6_, calc_stage_r_0__instr_operands__imm__5_, calc_stage_r_0__instr_operands__imm__4_, calc_stage_r_0__instr_operands__imm__3_, calc_stage_r_0__instr_operands__imm__2_, calc_stage_r_0__instr_operands__imm__1_, calc_stage_r_0__instr_operands__imm__0_ }),
    .exc_i({ exc_stage_r_0__poison_v_, exc_stage_r_0__roll_v_, exc_stage_r_0__illegal_instr_v_, exc_stage_r_0__tlb_miss_v_, exc_stage_r_0__load_fault_v_, exc_stage_r_0__store_fault_v_, exc_stage_r_0__cache_miss_v_ }),
    .mmu_cmd_o(mmu_cmd_o),
    .mmu_cmd_v_o(mmu_cmd_v_o),
    .mmu_cmd_ready_i(mmu_cmd_ready_i),
    .mmu_resp_i(mmu_resp_i),
    .mmu_resp_v_i(mmu_resp_v_i),
    .mmu_resp_ready_o(mmu_resp_ready_o),
    .result_o(mem_calc_result[127:64]),
    .cache_miss_o(exc_stage_n_3__cache_miss_v_)
  );


  bp_be_pipe_fp
  pipe_fp
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .decode_i({ calc_stage_r_0__decode__instr_v_, calc_stage_r_0__decode__fe_nop_v_, calc_stage_r_0__decode__be_nop_v_, calc_stage_r_0__decode__me_nop_v_, calc_stage_r_0__decode__pipe_comp_v_, calc_stage_r_0__decode__pipe_int_v_, calc_stage_r_0__decode__pipe_mul_v_, calc_stage_r_0__decode__pipe_mem_v_, calc_stage_r_0__decode__pipe_fp_v_, calc_stage_r_0__decode__irf_w_v_, calc_stage_r_0__decode__frf_w_v_, calc_stage_r_0__decode__mhartid_r_v_, calc_stage_r_0__decode__dcache_w_v_, calc_stage_r_0__decode__dcache_r_v_, calc_stage_r_0__decode__fp_not_int_v_, calc_stage_r_0__decode__ret_v_, calc_stage_r_0__decode__amo_v_, calc_stage_r_0__decode__jmp_v_, calc_stage_r_0__decode__br_v_, calc_stage_r_0__decode__opw_v_, calc_stage_r_0__decode__fu_op__fu_op__3_, calc_stage_r_0__decode__fu_op__fu_op__2_, calc_stage_r_0__decode__fu_op__fu_op__1_, calc_stage_r_0__decode__fu_op__fu_op__0_, calc_stage_r_0__decode__rs1_addr__4_, calc_stage_r_0__decode__rs1_addr__3_, calc_stage_r_0__decode__rs1_addr__2_, calc_stage_r_0__decode__rs1_addr__1_, calc_stage_r_0__decode__rs1_addr__0_, calc_stage_r_0__decode__rs2_addr__4_, calc_stage_r_0__decode__rs2_addr__3_, calc_stage_r_0__decode__rs2_addr__2_, calc_stage_r_0__decode__rs2_addr__1_, calc_stage_r_0__decode__rs2_addr__0_, calc_status_o[73:69], calc_stage_r_0__decode__src1_sel_, calc_stage_r_0__decode__src2_sel_, calc_stage_r_0__decode__baddr_sel_, calc_stage_r_0__decode__result_sel_ }),
    .rs1_i({ calc_stage_r_0__instr_operands__rs1__63_, calc_stage_r_0__instr_operands__rs1__62_, calc_stage_r_0__instr_operands__rs1__61_, calc_stage_r_0__instr_operands__rs1__60_, calc_stage_r_0__instr_operands__rs1__59_, calc_stage_r_0__instr_operands__rs1__58_, calc_stage_r_0__instr_operands__rs1__57_, calc_stage_r_0__instr_operands__rs1__56_, calc_stage_r_0__instr_operands__rs1__55_, calc_stage_r_0__instr_operands__rs1__54_, calc_stage_r_0__instr_operands__rs1__53_, calc_stage_r_0__instr_operands__rs1__52_, calc_stage_r_0__instr_operands__rs1__51_, calc_stage_r_0__instr_operands__rs1__50_, calc_stage_r_0__instr_operands__rs1__49_, calc_stage_r_0__instr_operands__rs1__48_, calc_stage_r_0__instr_operands__rs1__47_, calc_stage_r_0__instr_operands__rs1__46_, calc_stage_r_0__instr_operands__rs1__45_, calc_stage_r_0__instr_operands__rs1__44_, calc_stage_r_0__instr_operands__rs1__43_, calc_stage_r_0__instr_operands__rs1__42_, calc_stage_r_0__instr_operands__rs1__41_, calc_stage_r_0__instr_operands__rs1__40_, calc_stage_r_0__instr_operands__rs1__39_, calc_stage_r_0__instr_operands__rs1__38_, calc_stage_r_0__instr_operands__rs1__37_, calc_stage_r_0__instr_operands__rs1__36_, calc_stage_r_0__instr_operands__rs1__35_, calc_stage_r_0__instr_operands__rs1__34_, calc_stage_r_0__instr_operands__rs1__33_, calc_stage_r_0__instr_operands__rs1__32_, calc_stage_r_0__instr_operands__rs1__31_, calc_stage_r_0__instr_operands__rs1__30_, calc_stage_r_0__instr_operands__rs1__29_, calc_stage_r_0__instr_operands__rs1__28_, calc_stage_r_0__instr_operands__rs1__27_, calc_stage_r_0__instr_operands__rs1__26_, calc_stage_r_0__instr_operands__rs1__25_, calc_stage_r_0__instr_operands__rs1__24_, calc_stage_r_0__instr_operands__rs1__23_, calc_stage_r_0__instr_operands__rs1__22_, calc_stage_r_0__instr_operands__rs1__21_, calc_stage_r_0__instr_operands__rs1__20_, calc_stage_r_0__instr_operands__rs1__19_, calc_stage_r_0__instr_operands__rs1__18_, calc_stage_r_0__instr_operands__rs1__17_, calc_stage_r_0__instr_operands__rs1__16_, calc_stage_r_0__instr_operands__rs1__15_, calc_stage_r_0__instr_operands__rs1__14_, calc_stage_r_0__instr_operands__rs1__13_, calc_stage_r_0__instr_operands__rs1__12_, calc_stage_r_0__instr_operands__rs1__11_, calc_stage_r_0__instr_operands__rs1__10_, calc_stage_r_0__instr_operands__rs1__9_, calc_stage_r_0__instr_operands__rs1__8_, calc_stage_r_0__instr_operands__rs1__7_, calc_stage_r_0__instr_operands__rs1__6_, calc_stage_r_0__instr_operands__rs1__5_, calc_stage_r_0__instr_operands__rs1__4_, calc_stage_r_0__instr_operands__rs1__3_, calc_stage_r_0__instr_operands__rs1__2_, calc_stage_r_0__instr_operands__rs1__1_, calc_stage_r_0__instr_operands__rs1__0_ }),
    .rs2_i({ calc_stage_r_0__instr_operands__rs2__63_, calc_stage_r_0__instr_operands__rs2__62_, calc_stage_r_0__instr_operands__rs2__61_, calc_stage_r_0__instr_operands__rs2__60_, calc_stage_r_0__instr_operands__rs2__59_, calc_stage_r_0__instr_operands__rs2__58_, calc_stage_r_0__instr_operands__rs2__57_, calc_stage_r_0__instr_operands__rs2__56_, calc_stage_r_0__instr_operands__rs2__55_, calc_stage_r_0__instr_operands__rs2__54_, calc_stage_r_0__instr_operands__rs2__53_, calc_stage_r_0__instr_operands__rs2__52_, calc_stage_r_0__instr_operands__rs2__51_, calc_stage_r_0__instr_operands__rs2__50_, calc_stage_r_0__instr_operands__rs2__49_, calc_stage_r_0__instr_operands__rs2__48_, calc_stage_r_0__instr_operands__rs2__47_, calc_stage_r_0__instr_operands__rs2__46_, calc_stage_r_0__instr_operands__rs2__45_, calc_stage_r_0__instr_operands__rs2__44_, calc_stage_r_0__instr_operands__rs2__43_, calc_stage_r_0__instr_operands__rs2__42_, calc_stage_r_0__instr_operands__rs2__41_, calc_stage_r_0__instr_operands__rs2__40_, calc_stage_r_0__instr_operands__rs2__39_, calc_stage_r_0__instr_operands__rs2__38_, calc_stage_r_0__instr_operands__rs2__37_, calc_stage_r_0__instr_operands__rs2__36_, calc_stage_r_0__instr_operands__rs2__35_, calc_stage_r_0__instr_operands__rs2__34_, calc_stage_r_0__instr_operands__rs2__33_, calc_stage_r_0__instr_operands__rs2__32_, calc_stage_r_0__instr_operands__rs2__31_, calc_stage_r_0__instr_operands__rs2__30_, calc_stage_r_0__instr_operands__rs2__29_, calc_stage_r_0__instr_operands__rs2__28_, calc_stage_r_0__instr_operands__rs2__27_, calc_stage_r_0__instr_operands__rs2__26_, calc_stage_r_0__instr_operands__rs2__25_, calc_stage_r_0__instr_operands__rs2__24_, calc_stage_r_0__instr_operands__rs2__23_, calc_stage_r_0__instr_operands__rs2__22_, calc_stage_r_0__instr_operands__rs2__21_, calc_stage_r_0__instr_operands__rs2__20_, calc_stage_r_0__instr_operands__rs2__19_, calc_stage_r_0__instr_operands__rs2__18_, calc_stage_r_0__instr_operands__rs2__17_, calc_stage_r_0__instr_operands__rs2__16_, calc_stage_r_0__instr_operands__rs2__15_, calc_stage_r_0__instr_operands__rs2__14_, calc_stage_r_0__instr_operands__rs2__13_, calc_stage_r_0__instr_operands__rs2__12_, calc_stage_r_0__instr_operands__rs2__11_, calc_stage_r_0__instr_operands__rs2__10_, calc_stage_r_0__instr_operands__rs2__9_, calc_stage_r_0__instr_operands__rs2__8_, calc_stage_r_0__instr_operands__rs2__7_, calc_stage_r_0__instr_operands__rs2__6_, calc_stage_r_0__instr_operands__rs2__5_, calc_stage_r_0__instr_operands__rs2__4_, calc_stage_r_0__instr_operands__rs2__3_, calc_stage_r_0__instr_operands__rs2__2_, calc_stage_r_0__instr_operands__rs2__1_, calc_stage_r_0__instr_operands__rs2__0_ }),
    .exc_i({ exc_stage_r_0__poison_v_, exc_stage_r_0__roll_v_, exc_stage_r_0__illegal_instr_v_, exc_stage_r_0__tlb_miss_v_, exc_stage_r_0__load_fault_v_, exc_stage_r_0__store_fault_v_, exc_stage_r_0__cache_miss_v_ }),
    .result_o(fp_calc_result[127:64])
  );


  bsg_dff_width_p1890
  calc_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ calc_stage_r_3__instr_metadata__itag__7_, calc_stage_r_3__instr_metadata__itag__6_, calc_stage_r_3__instr_metadata__itag__5_, calc_stage_r_3__instr_metadata__itag__4_, calc_stage_r_3__instr_metadata__itag__3_, calc_stage_r_3__instr_metadata__itag__2_, calc_stage_r_3__instr_metadata__itag__1_, calc_stage_r_3__instr_metadata__itag__0_, calc_stage_r_3__instr_metadata__pc__63_, calc_stage_r_3__instr_metadata__pc__62_, calc_stage_r_3__instr_metadata__pc__61_, calc_stage_r_3__instr_metadata__pc__60_, calc_stage_r_3__instr_metadata__pc__59_, calc_stage_r_3__instr_metadata__pc__58_, calc_stage_r_3__instr_metadata__pc__57_, calc_stage_r_3__instr_metadata__pc__56_, calc_stage_r_3__instr_metadata__pc__55_, calc_stage_r_3__instr_metadata__pc__54_, calc_stage_r_3__instr_metadata__pc__53_, calc_stage_r_3__instr_metadata__pc__52_, calc_stage_r_3__instr_metadata__pc__51_, calc_stage_r_3__instr_metadata__pc__50_, calc_stage_r_3__instr_metadata__pc__49_, calc_stage_r_3__instr_metadata__pc__48_, calc_stage_r_3__instr_metadata__pc__47_, calc_stage_r_3__instr_metadata__pc__46_, calc_stage_r_3__instr_metadata__pc__45_, calc_stage_r_3__instr_metadata__pc__44_, calc_stage_r_3__instr_metadata__pc__43_, calc_stage_r_3__instr_metadata__pc__42_, calc_stage_r_3__instr_metadata__pc__41_, calc_stage_r_3__instr_metadata__pc__40_, calc_stage_r_3__instr_metadata__pc__39_, calc_stage_r_3__instr_metadata__pc__38_, calc_stage_r_3__instr_metadata__pc__37_, calc_stage_r_3__instr_metadata__pc__36_, calc_stage_r_3__instr_metadata__pc__35_, calc_stage_r_3__instr_metadata__pc__34_, calc_stage_r_3__instr_metadata__pc__33_, calc_stage_r_3__instr_metadata__pc__32_, calc_stage_r_3__instr_metadata__pc__31_, calc_stage_r_3__instr_metadata__pc__30_, calc_stage_r_3__instr_metadata__pc__29_, calc_stage_r_3__instr_metadata__pc__28_, calc_stage_r_3__instr_metadata__pc__27_, calc_stage_r_3__instr_metadata__pc__26_, calc_stage_r_3__instr_metadata__pc__25_, calc_stage_r_3__instr_metadata__pc__24_, calc_stage_r_3__instr_metadata__pc__23_, calc_stage_r_3__instr_metadata__pc__22_, calc_stage_r_3__instr_metadata__pc__21_, calc_stage_r_3__instr_metadata__pc__20_, calc_stage_r_3__instr_metadata__pc__19_, calc_stage_r_3__instr_metadata__pc__18_, calc_stage_r_3__instr_metadata__pc__17_, calc_stage_r_3__instr_metadata__pc__16_, calc_stage_r_3__instr_metadata__pc__15_, calc_stage_r_3__instr_metadata__pc__14_, calc_stage_r_3__instr_metadata__pc__13_, calc_stage_r_3__instr_metadata__pc__12_, calc_stage_r_3__instr_metadata__pc__11_, calc_stage_r_3__instr_metadata__pc__10_, calc_stage_r_3__instr_metadata__pc__9_, calc_stage_r_3__instr_metadata__pc__8_, calc_stage_r_3__instr_metadata__pc__7_, calc_stage_r_3__instr_metadata__pc__6_, calc_stage_r_3__instr_metadata__pc__5_, calc_stage_r_3__instr_metadata__pc__4_, calc_stage_r_3__instr_metadata__pc__3_, calc_stage_r_3__instr_metadata__pc__2_, calc_stage_r_3__instr_metadata__pc__1_, calc_stage_r_3__instr_metadata__pc__0_, calc_stage_r_3__instr_metadata__fe_exception_not_instr_, calc_stage_r_3__instr_metadata__fe_exception_code__1_, calc_stage_r_3__instr_metadata__fe_exception_code__0_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__35_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__34_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__33_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__32_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__31_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__30_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__29_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__28_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__27_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__26_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__25_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__24_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__23_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__22_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__21_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__20_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__19_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__18_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__17_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__16_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__15_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__14_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__13_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__12_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__11_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__10_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__9_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__8_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__7_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__6_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__5_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__4_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__3_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__2_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__1_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__0_, calc_stage_r_3__instr__31_, calc_stage_r_3__instr__30_, calc_stage_r_3__instr__29_, calc_stage_r_3__instr__28_, calc_stage_r_3__instr__27_, calc_stage_r_3__instr__26_, calc_stage_r_3__instr__25_, calc_stage_r_3__instr__24_, calc_stage_r_3__instr__23_, calc_stage_r_3__instr__22_, calc_stage_r_3__instr__21_, calc_stage_r_3__instr__20_, calc_stage_r_3__instr__19_, calc_stage_r_3__instr__18_, calc_stage_r_3__instr__17_, calc_stage_r_3__instr__16_, calc_stage_r_3__instr__15_, calc_stage_r_3__instr__14_, calc_stage_r_3__instr__13_, calc_stage_r_3__instr__12_, calc_stage_r_3__instr__11_, calc_stage_r_3__instr__10_, calc_stage_r_3__instr__9_, calc_stage_r_3__instr__8_, calc_stage_r_3__instr__7_, calc_stage_r_3__instr__6_, calc_stage_r_3__instr__5_, calc_stage_r_3__instr__4_, calc_stage_r_3__instr__3_, calc_stage_r_3__instr__2_, calc_stage_r_3__instr__1_, calc_stage_r_3__instr__0_, calc_stage_r_3__instr_operands__rs1__63_, calc_stage_r_3__instr_operands__rs1__62_, calc_stage_r_3__instr_operands__rs1__61_, calc_stage_r_3__instr_operands__rs1__60_, calc_stage_r_3__instr_operands__rs1__59_, calc_stage_r_3__instr_operands__rs1__58_, calc_stage_r_3__instr_operands__rs1__57_, calc_stage_r_3__instr_operands__rs1__56_, calc_stage_r_3__instr_operands__rs1__55_, calc_stage_r_3__instr_operands__rs1__54_, calc_stage_r_3__instr_operands__rs1__53_, calc_stage_r_3__instr_operands__rs1__52_, calc_stage_r_3__instr_operands__rs1__51_, calc_stage_r_3__instr_operands__rs1__50_, calc_stage_r_3__instr_operands__rs1__49_, calc_stage_r_3__instr_operands__rs1__48_, calc_stage_r_3__instr_operands__rs1__47_, calc_stage_r_3__instr_operands__rs1__46_, calc_stage_r_3__instr_operands__rs1__45_, calc_stage_r_3__instr_operands__rs1__44_, calc_stage_r_3__instr_operands__rs1__43_, calc_stage_r_3__instr_operands__rs1__42_, calc_stage_r_3__instr_operands__rs1__41_, calc_stage_r_3__instr_operands__rs1__40_, calc_stage_r_3__instr_operands__rs1__39_, calc_stage_r_3__instr_operands__rs1__38_, calc_stage_r_3__instr_operands__rs1__37_, calc_stage_r_3__instr_operands__rs1__36_, calc_stage_r_3__instr_operands__rs1__35_, calc_stage_r_3__instr_operands__rs1__34_, calc_stage_r_3__instr_operands__rs1__33_, calc_stage_r_3__instr_operands__rs1__32_, calc_stage_r_3__instr_operands__rs1__31_, calc_stage_r_3__instr_operands__rs1__30_, calc_stage_r_3__instr_operands__rs1__29_, calc_stage_r_3__instr_operands__rs1__28_, calc_stage_r_3__instr_operands__rs1__27_, calc_stage_r_3__instr_operands__rs1__26_, calc_stage_r_3__instr_operands__rs1__25_, calc_stage_r_3__instr_operands__rs1__24_, calc_stage_r_3__instr_operands__rs1__23_, calc_stage_r_3__instr_operands__rs1__22_, calc_stage_r_3__instr_operands__rs1__21_, calc_stage_r_3__instr_operands__rs1__20_, calc_stage_r_3__instr_operands__rs1__19_, calc_stage_r_3__instr_operands__rs1__18_, calc_stage_r_3__instr_operands__rs1__17_, calc_stage_r_3__instr_operands__rs1__16_, calc_stage_r_3__instr_operands__rs1__15_, calc_stage_r_3__instr_operands__rs1__14_, calc_stage_r_3__instr_operands__rs1__13_, calc_stage_r_3__instr_operands__rs1__12_, calc_stage_r_3__instr_operands__rs1__11_, calc_stage_r_3__instr_operands__rs1__10_, calc_stage_r_3__instr_operands__rs1__9_, calc_stage_r_3__instr_operands__rs1__8_, calc_stage_r_3__instr_operands__rs1__7_, calc_stage_r_3__instr_operands__rs1__6_, calc_stage_r_3__instr_operands__rs1__5_, calc_stage_r_3__instr_operands__rs1__4_, calc_stage_r_3__instr_operands__rs1__3_, calc_stage_r_3__instr_operands__rs1__2_, calc_stage_r_3__instr_operands__rs1__1_, calc_stage_r_3__instr_operands__rs1__0_, calc_stage_r_3__instr_operands__rs2__63_, calc_stage_r_3__instr_operands__rs2__62_, calc_stage_r_3__instr_operands__rs2__61_, calc_stage_r_3__instr_operands__rs2__60_, calc_stage_r_3__instr_operands__rs2__59_, calc_stage_r_3__instr_operands__rs2__58_, calc_stage_r_3__instr_operands__rs2__57_, calc_stage_r_3__instr_operands__rs2__56_, calc_stage_r_3__instr_operands__rs2__55_, calc_stage_r_3__instr_operands__rs2__54_, calc_stage_r_3__instr_operands__rs2__53_, calc_stage_r_3__instr_operands__rs2__52_, calc_stage_r_3__instr_operands__rs2__51_, calc_stage_r_3__instr_operands__rs2__50_, calc_stage_r_3__instr_operands__rs2__49_, calc_stage_r_3__instr_operands__rs2__48_, calc_stage_r_3__instr_operands__rs2__47_, calc_stage_r_3__instr_operands__rs2__46_, calc_stage_r_3__instr_operands__rs2__45_, calc_stage_r_3__instr_operands__rs2__44_, calc_stage_r_3__instr_operands__rs2__43_, calc_stage_r_3__instr_operands__rs2__42_, calc_stage_r_3__instr_operands__rs2__41_, calc_stage_r_3__instr_operands__rs2__40_, calc_stage_r_3__instr_operands__rs2__39_, calc_stage_r_3__instr_operands__rs2__38_, calc_stage_r_3__instr_operands__rs2__37_, calc_stage_r_3__instr_operands__rs2__36_, calc_stage_r_3__instr_operands__rs2__35_, calc_stage_r_3__instr_operands__rs2__34_, calc_stage_r_3__instr_operands__rs2__33_, calc_stage_r_3__instr_operands__rs2__32_, calc_stage_r_3__instr_operands__rs2__31_, calc_stage_r_3__instr_operands__rs2__30_, calc_stage_r_3__instr_operands__rs2__29_, calc_stage_r_3__instr_operands__rs2__28_, calc_stage_r_3__instr_operands__rs2__27_, calc_stage_r_3__instr_operands__rs2__26_, calc_stage_r_3__instr_operands__rs2__25_, calc_stage_r_3__instr_operands__rs2__24_, calc_stage_r_3__instr_operands__rs2__23_, calc_stage_r_3__instr_operands__rs2__22_, calc_stage_r_3__instr_operands__rs2__21_, calc_stage_r_3__instr_operands__rs2__20_, calc_stage_r_3__instr_operands__rs2__19_, calc_stage_r_3__instr_operands__rs2__18_, calc_stage_r_3__instr_operands__rs2__17_, calc_stage_r_3__instr_operands__rs2__16_, calc_stage_r_3__instr_operands__rs2__15_, calc_stage_r_3__instr_operands__rs2__14_, calc_stage_r_3__instr_operands__rs2__13_, calc_stage_r_3__instr_operands__rs2__12_, calc_stage_r_3__instr_operands__rs2__11_, calc_stage_r_3__instr_operands__rs2__10_, calc_stage_r_3__instr_operands__rs2__9_, calc_stage_r_3__instr_operands__rs2__8_, calc_stage_r_3__instr_operands__rs2__7_, calc_stage_r_3__instr_operands__rs2__6_, calc_stage_r_3__instr_operands__rs2__5_, calc_stage_r_3__instr_operands__rs2__4_, calc_stage_r_3__instr_operands__rs2__3_, calc_stage_r_3__instr_operands__rs2__2_, calc_stage_r_3__instr_operands__rs2__1_, calc_stage_r_3__instr_operands__rs2__0_, calc_stage_r_3__instr_operands__imm__63_, calc_stage_r_3__instr_operands__imm__62_, calc_stage_r_3__instr_operands__imm__61_, calc_stage_r_3__instr_operands__imm__60_, calc_stage_r_3__instr_operands__imm__59_, calc_stage_r_3__instr_operands__imm__58_, calc_stage_r_3__instr_operands__imm__57_, calc_stage_r_3__instr_operands__imm__56_, calc_stage_r_3__instr_operands__imm__55_, calc_stage_r_3__instr_operands__imm__54_, calc_stage_r_3__instr_operands__imm__53_, calc_stage_r_3__instr_operands__imm__52_, calc_stage_r_3__instr_operands__imm__51_, calc_stage_r_3__instr_operands__imm__50_, calc_stage_r_3__instr_operands__imm__49_, calc_stage_r_3__instr_operands__imm__48_, calc_stage_r_3__instr_operands__imm__47_, calc_stage_r_3__instr_operands__imm__46_, calc_stage_r_3__instr_operands__imm__45_, calc_stage_r_3__instr_operands__imm__44_, calc_stage_r_3__instr_operands__imm__43_, calc_stage_r_3__instr_operands__imm__42_, calc_stage_r_3__instr_operands__imm__41_, calc_stage_r_3__instr_operands__imm__40_, calc_stage_r_3__instr_operands__imm__39_, calc_stage_r_3__instr_operands__imm__38_, calc_stage_r_3__instr_operands__imm__37_, calc_stage_r_3__instr_operands__imm__36_, calc_stage_r_3__instr_operands__imm__35_, calc_stage_r_3__instr_operands__imm__34_, calc_stage_r_3__instr_operands__imm__33_, calc_stage_r_3__instr_operands__imm__32_, calc_stage_r_3__instr_operands__imm__31_, calc_stage_r_3__instr_operands__imm__30_, calc_stage_r_3__instr_operands__imm__29_, calc_stage_r_3__instr_operands__imm__28_, calc_stage_r_3__instr_operands__imm__27_, calc_stage_r_3__instr_operands__imm__26_, calc_stage_r_3__instr_operands__imm__25_, calc_stage_r_3__instr_operands__imm__24_, calc_stage_r_3__instr_operands__imm__23_, calc_stage_r_3__instr_operands__imm__22_, calc_stage_r_3__instr_operands__imm__21_, calc_stage_r_3__instr_operands__imm__20_, calc_stage_r_3__instr_operands__imm__19_, calc_stage_r_3__instr_operands__imm__18_, calc_stage_r_3__instr_operands__imm__17_, calc_stage_r_3__instr_operands__imm__16_, calc_stage_r_3__instr_operands__imm__15_, calc_stage_r_3__instr_operands__imm__14_, calc_stage_r_3__instr_operands__imm__13_, calc_stage_r_3__instr_operands__imm__12_, calc_stage_r_3__instr_operands__imm__11_, calc_stage_r_3__instr_operands__imm__10_, calc_stage_r_3__instr_operands__imm__9_, calc_stage_r_3__instr_operands__imm__8_, calc_stage_r_3__instr_operands__imm__7_, calc_stage_r_3__instr_operands__imm__6_, calc_stage_r_3__instr_operands__imm__5_, calc_stage_r_3__instr_operands__imm__4_, calc_stage_r_3__instr_operands__imm__3_, calc_stage_r_3__instr_operands__imm__2_, calc_stage_r_3__instr_operands__imm__1_, calc_stage_r_3__instr_operands__imm__0_, calc_stage_r_3__decode__instr_v_, calc_stage_r_3__decode__fe_nop_v_, calc_stage_r_3__decode__be_nop_v_, calc_stage_r_3__decode__me_nop_v_, calc_stage_r_3__decode__pipe_comp_v_, calc_stage_r_3__decode__pipe_int_v_, calc_stage_r_3__decode__pipe_mul_v_, calc_stage_r_3__decode__pipe_mem_v_, calc_stage_r_3__decode__pipe_fp_v_, calc_stage_r_3__decode__irf_w_v_, calc_stage_r_3__decode__frf_w_v_, calc_stage_r_3__decode__mhartid_r_v_, calc_stage_r_3__decode__dcache_w_v_, calc_stage_r_3__decode__dcache_r_v_, calc_stage_r_3__decode__fp_not_int_v_, calc_stage_r_3__decode__ret_v_, calc_stage_r_3__decode__amo_v_, calc_stage_r_3__decode__jmp_v_, calc_stage_r_3__decode__br_v_, calc_stage_r_3__decode__opw_v_, calc_stage_r_3__decode__fu_op__fu_op__3_, calc_stage_r_3__decode__fu_op__fu_op__2_, calc_stage_r_3__decode__fu_op__fu_op__1_, calc_stage_r_3__decode__fu_op__fu_op__0_, calc_stage_r_3__decode__rs1_addr__4_, calc_stage_r_3__decode__rs1_addr__3_, calc_stage_r_3__decode__rs1_addr__2_, calc_stage_r_3__decode__rs1_addr__1_, calc_stage_r_3__decode__rs1_addr__0_, calc_stage_r_3__decode__rs2_addr__4_, calc_stage_r_3__decode__rs2_addr__3_, calc_stage_r_3__decode__rs2_addr__2_, calc_stage_r_3__decode__rs2_addr__1_, calc_stage_r_3__decode__rs2_addr__0_, calc_status_o[103:99], calc_stage_r_3__decode__src1_sel_, calc_stage_r_3__decode__src2_sel_, calc_stage_r_3__decode__baddr_sel_, calc_stage_r_3__decode__result_sel_, calc_stage_r_2__instr_metadata__itag__7_, calc_stage_r_2__instr_metadata__itag__6_, calc_stage_r_2__instr_metadata__itag__5_, calc_stage_r_2__instr_metadata__itag__4_, calc_stage_r_2__instr_metadata__itag__3_, calc_stage_r_2__instr_metadata__itag__2_, calc_stage_r_2__instr_metadata__itag__1_, calc_stage_r_2__instr_metadata__itag__0_, calc_status_o[67:4], calc_stage_r_2__instr_metadata__fe_exception_not_instr_, calc_stage_r_2__instr_metadata__fe_exception_code__1_, calc_stage_r_2__instr_metadata__fe_exception_code__0_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__35_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__34_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__33_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__32_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__31_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__30_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__29_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__28_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__27_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__26_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__25_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__24_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__23_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__22_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__21_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__20_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__19_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__18_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__17_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__16_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__15_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__14_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__13_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__12_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__11_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__10_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__9_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__8_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__7_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__6_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__5_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__4_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__3_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__2_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__1_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__0_, calc_stage_r_2__instr__31_, calc_stage_r_2__instr__30_, calc_stage_r_2__instr__29_, calc_stage_r_2__instr__28_, calc_stage_r_2__instr__27_, calc_stage_r_2__instr__26_, calc_stage_r_2__instr__25_, calc_stage_r_2__instr__24_, calc_stage_r_2__instr__23_, calc_stage_r_2__instr__22_, calc_stage_r_2__instr__21_, calc_stage_r_2__instr__20_, calc_stage_r_2__instr__19_, calc_stage_r_2__instr__18_, calc_stage_r_2__instr__17_, calc_stage_r_2__instr__16_, calc_stage_r_2__instr__15_, calc_stage_r_2__instr__14_, calc_stage_r_2__instr__13_, calc_stage_r_2__instr__12_, calc_stage_r_2__instr__11_, calc_stage_r_2__instr__10_, calc_stage_r_2__instr__9_, calc_stage_r_2__instr__8_, calc_stage_r_2__instr__7_, calc_stage_r_2__instr__6_, calc_stage_r_2__instr__5_, calc_stage_r_2__instr__4_, calc_stage_r_2__instr__3_, calc_stage_r_2__instr__2_, calc_stage_r_2__instr__1_, calc_stage_r_2__instr__0_, calc_stage_r_2__instr_operands__rs1__63_, calc_stage_r_2__instr_operands__rs1__62_, calc_stage_r_2__instr_operands__rs1__61_, calc_stage_r_2__instr_operands__rs1__60_, calc_stage_r_2__instr_operands__rs1__59_, calc_stage_r_2__instr_operands__rs1__58_, calc_stage_r_2__instr_operands__rs1__57_, calc_stage_r_2__instr_operands__rs1__56_, calc_stage_r_2__instr_operands__rs1__55_, calc_stage_r_2__instr_operands__rs1__54_, calc_stage_r_2__instr_operands__rs1__53_, calc_stage_r_2__instr_operands__rs1__52_, calc_stage_r_2__instr_operands__rs1__51_, calc_stage_r_2__instr_operands__rs1__50_, calc_stage_r_2__instr_operands__rs1__49_, calc_stage_r_2__instr_operands__rs1__48_, calc_stage_r_2__instr_operands__rs1__47_, calc_stage_r_2__instr_operands__rs1__46_, calc_stage_r_2__instr_operands__rs1__45_, calc_stage_r_2__instr_operands__rs1__44_, calc_stage_r_2__instr_operands__rs1__43_, calc_stage_r_2__instr_operands__rs1__42_, calc_stage_r_2__instr_operands__rs1__41_, calc_stage_r_2__instr_operands__rs1__40_, calc_stage_r_2__instr_operands__rs1__39_, calc_stage_r_2__instr_operands__rs1__38_, calc_stage_r_2__instr_operands__rs1__37_, calc_stage_r_2__instr_operands__rs1__36_, calc_stage_r_2__instr_operands__rs1__35_, calc_stage_r_2__instr_operands__rs1__34_, calc_stage_r_2__instr_operands__rs1__33_, calc_stage_r_2__instr_operands__rs1__32_, calc_stage_r_2__instr_operands__rs1__31_, calc_stage_r_2__instr_operands__rs1__30_, calc_stage_r_2__instr_operands__rs1__29_, calc_stage_r_2__instr_operands__rs1__28_, calc_stage_r_2__instr_operands__rs1__27_, calc_stage_r_2__instr_operands__rs1__26_, calc_stage_r_2__instr_operands__rs1__25_, calc_stage_r_2__instr_operands__rs1__24_, calc_stage_r_2__instr_operands__rs1__23_, calc_stage_r_2__instr_operands__rs1__22_, calc_stage_r_2__instr_operands__rs1__21_, calc_stage_r_2__instr_operands__rs1__20_, calc_stage_r_2__instr_operands__rs1__19_, calc_stage_r_2__instr_operands__rs1__18_, calc_stage_r_2__instr_operands__rs1__17_, calc_stage_r_2__instr_operands__rs1__16_, calc_stage_r_2__instr_operands__rs1__15_, calc_stage_r_2__instr_operands__rs1__14_, calc_stage_r_2__instr_operands__rs1__13_, calc_stage_r_2__instr_operands__rs1__12_, calc_stage_r_2__instr_operands__rs1__11_, calc_stage_r_2__instr_operands__rs1__10_, calc_stage_r_2__instr_operands__rs1__9_, calc_stage_r_2__instr_operands__rs1__8_, calc_stage_r_2__instr_operands__rs1__7_, calc_stage_r_2__instr_operands__rs1__6_, calc_stage_r_2__instr_operands__rs1__5_, calc_stage_r_2__instr_operands__rs1__4_, calc_stage_r_2__instr_operands__rs1__3_, calc_stage_r_2__instr_operands__rs1__2_, calc_stage_r_2__instr_operands__rs1__1_, calc_stage_r_2__instr_operands__rs1__0_, calc_stage_r_2__instr_operands__rs2__63_, calc_stage_r_2__instr_operands__rs2__62_, calc_stage_r_2__instr_operands__rs2__61_, calc_stage_r_2__instr_operands__rs2__60_, calc_stage_r_2__instr_operands__rs2__59_, calc_stage_r_2__instr_operands__rs2__58_, calc_stage_r_2__instr_operands__rs2__57_, calc_stage_r_2__instr_operands__rs2__56_, calc_stage_r_2__instr_operands__rs2__55_, calc_stage_r_2__instr_operands__rs2__54_, calc_stage_r_2__instr_operands__rs2__53_, calc_stage_r_2__instr_operands__rs2__52_, calc_stage_r_2__instr_operands__rs2__51_, calc_stage_r_2__instr_operands__rs2__50_, calc_stage_r_2__instr_operands__rs2__49_, calc_stage_r_2__instr_operands__rs2__48_, calc_stage_r_2__instr_operands__rs2__47_, calc_stage_r_2__instr_operands__rs2__46_, calc_stage_r_2__instr_operands__rs2__45_, calc_stage_r_2__instr_operands__rs2__44_, calc_stage_r_2__instr_operands__rs2__43_, calc_stage_r_2__instr_operands__rs2__42_, calc_stage_r_2__instr_operands__rs2__41_, calc_stage_r_2__instr_operands__rs2__40_, calc_stage_r_2__instr_operands__rs2__39_, calc_stage_r_2__instr_operands__rs2__38_, calc_stage_r_2__instr_operands__rs2__37_, calc_stage_r_2__instr_operands__rs2__36_, calc_stage_r_2__instr_operands__rs2__35_, calc_stage_r_2__instr_operands__rs2__34_, calc_stage_r_2__instr_operands__rs2__33_, calc_stage_r_2__instr_operands__rs2__32_, calc_stage_r_2__instr_operands__rs2__31_, calc_stage_r_2__instr_operands__rs2__30_, calc_stage_r_2__instr_operands__rs2__29_, calc_stage_r_2__instr_operands__rs2__28_, calc_stage_r_2__instr_operands__rs2__27_, calc_stage_r_2__instr_operands__rs2__26_, calc_stage_r_2__instr_operands__rs2__25_, calc_stage_r_2__instr_operands__rs2__24_, calc_stage_r_2__instr_operands__rs2__23_, calc_stage_r_2__instr_operands__rs2__22_, calc_stage_r_2__instr_operands__rs2__21_, calc_stage_r_2__instr_operands__rs2__20_, calc_stage_r_2__instr_operands__rs2__19_, calc_stage_r_2__instr_operands__rs2__18_, calc_stage_r_2__instr_operands__rs2__17_, calc_stage_r_2__instr_operands__rs2__16_, calc_stage_r_2__instr_operands__rs2__15_, calc_stage_r_2__instr_operands__rs2__14_, calc_stage_r_2__instr_operands__rs2__13_, calc_stage_r_2__instr_operands__rs2__12_, calc_stage_r_2__instr_operands__rs2__11_, calc_stage_r_2__instr_operands__rs2__10_, calc_stage_r_2__instr_operands__rs2__9_, calc_stage_r_2__instr_operands__rs2__8_, calc_stage_r_2__instr_operands__rs2__7_, calc_stage_r_2__instr_operands__rs2__6_, calc_stage_r_2__instr_operands__rs2__5_, calc_stage_r_2__instr_operands__rs2__4_, calc_stage_r_2__instr_operands__rs2__3_, calc_stage_r_2__instr_operands__rs2__2_, calc_stage_r_2__instr_operands__rs2__1_, calc_stage_r_2__instr_operands__rs2__0_, calc_stage_r_2__instr_operands__imm__63_, calc_stage_r_2__instr_operands__imm__62_, calc_stage_r_2__instr_operands__imm__61_, calc_stage_r_2__instr_operands__imm__60_, calc_stage_r_2__instr_operands__imm__59_, calc_stage_r_2__instr_operands__imm__58_, calc_stage_r_2__instr_operands__imm__57_, calc_stage_r_2__instr_operands__imm__56_, calc_stage_r_2__instr_operands__imm__55_, calc_stage_r_2__instr_operands__imm__54_, calc_stage_r_2__instr_operands__imm__53_, calc_stage_r_2__instr_operands__imm__52_, calc_stage_r_2__instr_operands__imm__51_, calc_stage_r_2__instr_operands__imm__50_, calc_stage_r_2__instr_operands__imm__49_, calc_stage_r_2__instr_operands__imm__48_, calc_stage_r_2__instr_operands__imm__47_, calc_stage_r_2__instr_operands__imm__46_, calc_stage_r_2__instr_operands__imm__45_, calc_stage_r_2__instr_operands__imm__44_, calc_stage_r_2__instr_operands__imm__43_, calc_stage_r_2__instr_operands__imm__42_, calc_stage_r_2__instr_operands__imm__41_, calc_stage_r_2__instr_operands__imm__40_, calc_stage_r_2__instr_operands__imm__39_, calc_stage_r_2__instr_operands__imm__38_, calc_stage_r_2__instr_operands__imm__37_, calc_stage_r_2__instr_operands__imm__36_, calc_stage_r_2__instr_operands__imm__35_, calc_stage_r_2__instr_operands__imm__34_, calc_stage_r_2__instr_operands__imm__33_, calc_stage_r_2__instr_operands__imm__32_, calc_stage_r_2__instr_operands__imm__31_, calc_stage_r_2__instr_operands__imm__30_, calc_stage_r_2__instr_operands__imm__29_, calc_stage_r_2__instr_operands__imm__28_, calc_stage_r_2__instr_operands__imm__27_, calc_stage_r_2__instr_operands__imm__26_, calc_stage_r_2__instr_operands__imm__25_, calc_stage_r_2__instr_operands__imm__24_, calc_stage_r_2__instr_operands__imm__23_, calc_stage_r_2__instr_operands__imm__22_, calc_stage_r_2__instr_operands__imm__21_, calc_stage_r_2__instr_operands__imm__20_, calc_stage_r_2__instr_operands__imm__19_, calc_stage_r_2__instr_operands__imm__18_, calc_stage_r_2__instr_operands__imm__17_, calc_stage_r_2__instr_operands__imm__16_, calc_stage_r_2__instr_operands__imm__15_, calc_stage_r_2__instr_operands__imm__14_, calc_stage_r_2__instr_operands__imm__13_, calc_stage_r_2__instr_operands__imm__12_, calc_stage_r_2__instr_operands__imm__11_, calc_stage_r_2__instr_operands__imm__10_, calc_stage_r_2__instr_operands__imm__9_, calc_stage_r_2__instr_operands__imm__8_, calc_stage_r_2__instr_operands__imm__7_, calc_stage_r_2__instr_operands__imm__6_, calc_stage_r_2__instr_operands__imm__5_, calc_stage_r_2__instr_operands__imm__4_, calc_stage_r_2__instr_operands__imm__3_, calc_stage_r_2__instr_operands__imm__2_, calc_stage_r_2__instr_operands__imm__1_, calc_stage_r_2__instr_operands__imm__0_, calc_stage_r_2__decode__instr_v_, calc_stage_r_2__decode__fe_nop_v_, calc_stage_r_2__decode__be_nop_v_, calc_stage_r_2__decode__me_nop_v_, calc_stage_r_2__decode__pipe_comp_v_, calc_stage_r_2__decode__pipe_int_v_, calc_stage_r_2__decode__pipe_mul_v_, calc_stage_r_2__decode__pipe_mem_v_, calc_stage_r_2__decode__pipe_fp_v_, calc_stage_r_2__decode__irf_w_v_, calc_stage_r_2__decode__frf_w_v_, calc_stage_r_2__decode__mhartid_r_v_, calc_stage_r_2__decode__dcache_w_v_, calc_stage_r_2__decode__dcache_r_v_, calc_stage_r_2__decode__fp_not_int_v_, calc_status_o[1:1], calc_stage_r_2__decode__amo_v_, calc_stage_r_2__decode__jmp_v_, calc_stage_r_2__decode__br_v_, calc_stage_r_2__decode__opw_v_, calc_stage_r_2__decode__fu_op__fu_op__3_, calc_stage_r_2__decode__fu_op__fu_op__2_, calc_stage_r_2__decode__fu_op__fu_op__1_, calc_stage_r_2__decode__fu_op__fu_op__0_, calc_stage_r_2__decode__rs1_addr__4_, calc_stage_r_2__decode__rs1_addr__3_, calc_stage_r_2__decode__rs1_addr__2_, calc_stage_r_2__decode__rs1_addr__1_, calc_stage_r_2__decode__rs1_addr__0_, calc_stage_r_2__decode__rs2_addr__4_, calc_stage_r_2__decode__rs2_addr__3_, calc_stage_r_2__decode__rs2_addr__2_, calc_stage_r_2__decode__rs2_addr__1_, calc_stage_r_2__decode__rs2_addr__0_, calc_status_o[93:89], calc_stage_r_2__decode__src1_sel_, calc_stage_r_2__decode__src2_sel_, calc_stage_r_2__decode__baddr_sel_, calc_stage_r_2__decode__result_sel_, calc_stage_r_1__instr_metadata__itag__7_, calc_stage_r_1__instr_metadata__itag__6_, calc_stage_r_1__instr_metadata__itag__5_, calc_stage_r_1__instr_metadata__itag__4_, calc_stage_r_1__instr_metadata__itag__3_, calc_stage_r_1__instr_metadata__itag__2_, calc_stage_r_1__instr_metadata__itag__1_, calc_stage_r_1__instr_metadata__itag__0_, calc_stage_r_1__instr_metadata__pc__63_, calc_stage_r_1__instr_metadata__pc__62_, calc_stage_r_1__instr_metadata__pc__61_, calc_stage_r_1__instr_metadata__pc__60_, calc_stage_r_1__instr_metadata__pc__59_, calc_stage_r_1__instr_metadata__pc__58_, calc_stage_r_1__instr_metadata__pc__57_, calc_stage_r_1__instr_metadata__pc__56_, calc_stage_r_1__instr_metadata__pc__55_, calc_stage_r_1__instr_metadata__pc__54_, calc_stage_r_1__instr_metadata__pc__53_, calc_stage_r_1__instr_metadata__pc__52_, calc_stage_r_1__instr_metadata__pc__51_, calc_stage_r_1__instr_metadata__pc__50_, calc_stage_r_1__instr_metadata__pc__49_, calc_stage_r_1__instr_metadata__pc__48_, calc_stage_r_1__instr_metadata__pc__47_, calc_stage_r_1__instr_metadata__pc__46_, calc_stage_r_1__instr_metadata__pc__45_, calc_stage_r_1__instr_metadata__pc__44_, calc_stage_r_1__instr_metadata__pc__43_, calc_stage_r_1__instr_metadata__pc__42_, calc_stage_r_1__instr_metadata__pc__41_, calc_stage_r_1__instr_metadata__pc__40_, calc_stage_r_1__instr_metadata__pc__39_, calc_stage_r_1__instr_metadata__pc__38_, calc_stage_r_1__instr_metadata__pc__37_, calc_stage_r_1__instr_metadata__pc__36_, calc_stage_r_1__instr_metadata__pc__35_, calc_stage_r_1__instr_metadata__pc__34_, calc_stage_r_1__instr_metadata__pc__33_, calc_stage_r_1__instr_metadata__pc__32_, calc_stage_r_1__instr_metadata__pc__31_, calc_stage_r_1__instr_metadata__pc__30_, calc_stage_r_1__instr_metadata__pc__29_, calc_stage_r_1__instr_metadata__pc__28_, calc_stage_r_1__instr_metadata__pc__27_, calc_stage_r_1__instr_metadata__pc__26_, calc_stage_r_1__instr_metadata__pc__25_, calc_stage_r_1__instr_metadata__pc__24_, calc_stage_r_1__instr_metadata__pc__23_, calc_stage_r_1__instr_metadata__pc__22_, calc_stage_r_1__instr_metadata__pc__21_, calc_stage_r_1__instr_metadata__pc__20_, calc_stage_r_1__instr_metadata__pc__19_, calc_stage_r_1__instr_metadata__pc__18_, calc_stage_r_1__instr_metadata__pc__17_, calc_stage_r_1__instr_metadata__pc__16_, calc_stage_r_1__instr_metadata__pc__15_, calc_stage_r_1__instr_metadata__pc__14_, calc_stage_r_1__instr_metadata__pc__13_, calc_stage_r_1__instr_metadata__pc__12_, calc_stage_r_1__instr_metadata__pc__11_, calc_stage_r_1__instr_metadata__pc__10_, calc_stage_r_1__instr_metadata__pc__9_, calc_stage_r_1__instr_metadata__pc__8_, calc_stage_r_1__instr_metadata__pc__7_, calc_stage_r_1__instr_metadata__pc__6_, calc_stage_r_1__instr_metadata__pc__5_, calc_stage_r_1__instr_metadata__pc__4_, calc_stage_r_1__instr_metadata__pc__3_, calc_stage_r_1__instr_metadata__pc__2_, calc_stage_r_1__instr_metadata__pc__1_, calc_stage_r_1__instr_metadata__pc__0_, calc_stage_r_1__instr_metadata__fe_exception_not_instr_, calc_stage_r_1__instr_metadata__fe_exception_code__1_, calc_stage_r_1__instr_metadata__fe_exception_code__0_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__35_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__34_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__33_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__32_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__31_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__30_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__29_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__28_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__27_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__26_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__25_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__24_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__23_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__22_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__21_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__20_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__19_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__18_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__17_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__16_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__15_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__14_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__13_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__12_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__11_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__10_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__9_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__8_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__7_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__6_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__5_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__4_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__3_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__2_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__1_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__0_, calc_stage_r_1__instr__31_, calc_stage_r_1__instr__30_, calc_stage_r_1__instr__29_, calc_stage_r_1__instr__28_, calc_stage_r_1__instr__27_, calc_stage_r_1__instr__26_, calc_stage_r_1__instr__25_, calc_stage_r_1__instr__24_, calc_stage_r_1__instr__23_, calc_stage_r_1__instr__22_, calc_stage_r_1__instr__21_, calc_stage_r_1__instr__20_, calc_stage_r_1__instr__19_, calc_stage_r_1__instr__18_, calc_stage_r_1__instr__17_, calc_stage_r_1__instr__16_, calc_stage_r_1__instr__15_, calc_stage_r_1__instr__14_, calc_stage_r_1__instr__13_, calc_stage_r_1__instr__12_, calc_stage_r_1__instr__11_, calc_stage_r_1__instr__10_, calc_stage_r_1__instr__9_, calc_stage_r_1__instr__8_, calc_stage_r_1__instr__7_, calc_stage_r_1__instr__6_, calc_stage_r_1__instr__5_, calc_stage_r_1__instr__4_, calc_stage_r_1__instr__3_, calc_stage_r_1__instr__2_, calc_stage_r_1__instr__1_, calc_stage_r_1__instr__0_, calc_stage_r_1__instr_operands__rs1__63_, calc_stage_r_1__instr_operands__rs1__62_, calc_stage_r_1__instr_operands__rs1__61_, calc_stage_r_1__instr_operands__rs1__60_, calc_stage_r_1__instr_operands__rs1__59_, calc_stage_r_1__instr_operands__rs1__58_, calc_stage_r_1__instr_operands__rs1__57_, calc_stage_r_1__instr_operands__rs1__56_, calc_stage_r_1__instr_operands__rs1__55_, calc_stage_r_1__instr_operands__rs1__54_, calc_stage_r_1__instr_operands__rs1__53_, calc_stage_r_1__instr_operands__rs1__52_, calc_stage_r_1__instr_operands__rs1__51_, calc_stage_r_1__instr_operands__rs1__50_, calc_stage_r_1__instr_operands__rs1__49_, calc_stage_r_1__instr_operands__rs1__48_, calc_stage_r_1__instr_operands__rs1__47_, calc_stage_r_1__instr_operands__rs1__46_, calc_stage_r_1__instr_operands__rs1__45_, calc_stage_r_1__instr_operands__rs1__44_, calc_stage_r_1__instr_operands__rs1__43_, calc_stage_r_1__instr_operands__rs1__42_, calc_stage_r_1__instr_operands__rs1__41_, calc_stage_r_1__instr_operands__rs1__40_, calc_stage_r_1__instr_operands__rs1__39_, calc_stage_r_1__instr_operands__rs1__38_, calc_stage_r_1__instr_operands__rs1__37_, calc_stage_r_1__instr_operands__rs1__36_, calc_stage_r_1__instr_operands__rs1__35_, calc_stage_r_1__instr_operands__rs1__34_, calc_stage_r_1__instr_operands__rs1__33_, calc_stage_r_1__instr_operands__rs1__32_, calc_stage_r_1__instr_operands__rs1__31_, calc_stage_r_1__instr_operands__rs1__30_, calc_stage_r_1__instr_operands__rs1__29_, calc_stage_r_1__instr_operands__rs1__28_, calc_stage_r_1__instr_operands__rs1__27_, calc_stage_r_1__instr_operands__rs1__26_, calc_stage_r_1__instr_operands__rs1__25_, calc_stage_r_1__instr_operands__rs1__24_, calc_stage_r_1__instr_operands__rs1__23_, calc_stage_r_1__instr_operands__rs1__22_, calc_stage_r_1__instr_operands__rs1__21_, calc_stage_r_1__instr_operands__rs1__20_, calc_stage_r_1__instr_operands__rs1__19_, calc_stage_r_1__instr_operands__rs1__18_, calc_stage_r_1__instr_operands__rs1__17_, calc_stage_r_1__instr_operands__rs1__16_, calc_stage_r_1__instr_operands__rs1__15_, calc_stage_r_1__instr_operands__rs1__14_, calc_stage_r_1__instr_operands__rs1__13_, calc_stage_r_1__instr_operands__rs1__12_, calc_stage_r_1__instr_operands__rs1__11_, calc_stage_r_1__instr_operands__rs1__10_, calc_stage_r_1__instr_operands__rs1__9_, calc_stage_r_1__instr_operands__rs1__8_, calc_stage_r_1__instr_operands__rs1__7_, calc_stage_r_1__instr_operands__rs1__6_, calc_stage_r_1__instr_operands__rs1__5_, calc_stage_r_1__instr_operands__rs1__4_, calc_stage_r_1__instr_operands__rs1__3_, calc_stage_r_1__instr_operands__rs1__2_, calc_stage_r_1__instr_operands__rs1__1_, calc_stage_r_1__instr_operands__rs1__0_, calc_stage_r_1__instr_operands__rs2__63_, calc_stage_r_1__instr_operands__rs2__62_, calc_stage_r_1__instr_operands__rs2__61_, calc_stage_r_1__instr_operands__rs2__60_, calc_stage_r_1__instr_operands__rs2__59_, calc_stage_r_1__instr_operands__rs2__58_, calc_stage_r_1__instr_operands__rs2__57_, calc_stage_r_1__instr_operands__rs2__56_, calc_stage_r_1__instr_operands__rs2__55_, calc_stage_r_1__instr_operands__rs2__54_, calc_stage_r_1__instr_operands__rs2__53_, calc_stage_r_1__instr_operands__rs2__52_, calc_stage_r_1__instr_operands__rs2__51_, calc_stage_r_1__instr_operands__rs2__50_, calc_stage_r_1__instr_operands__rs2__49_, calc_stage_r_1__instr_operands__rs2__48_, calc_stage_r_1__instr_operands__rs2__47_, calc_stage_r_1__instr_operands__rs2__46_, calc_stage_r_1__instr_operands__rs2__45_, calc_stage_r_1__instr_operands__rs2__44_, calc_stage_r_1__instr_operands__rs2__43_, calc_stage_r_1__instr_operands__rs2__42_, calc_stage_r_1__instr_operands__rs2__41_, calc_stage_r_1__instr_operands__rs2__40_, calc_stage_r_1__instr_operands__rs2__39_, calc_stage_r_1__instr_operands__rs2__38_, calc_stage_r_1__instr_operands__rs2__37_, calc_stage_r_1__instr_operands__rs2__36_, calc_stage_r_1__instr_operands__rs2__35_, calc_stage_r_1__instr_operands__rs2__34_, calc_stage_r_1__instr_operands__rs2__33_, calc_stage_r_1__instr_operands__rs2__32_, calc_stage_r_1__instr_operands__rs2__31_, calc_stage_r_1__instr_operands__rs2__30_, calc_stage_r_1__instr_operands__rs2__29_, calc_stage_r_1__instr_operands__rs2__28_, calc_stage_r_1__instr_operands__rs2__27_, calc_stage_r_1__instr_operands__rs2__26_, calc_stage_r_1__instr_operands__rs2__25_, calc_stage_r_1__instr_operands__rs2__24_, calc_stage_r_1__instr_operands__rs2__23_, calc_stage_r_1__instr_operands__rs2__22_, calc_stage_r_1__instr_operands__rs2__21_, calc_stage_r_1__instr_operands__rs2__20_, calc_stage_r_1__instr_operands__rs2__19_, calc_stage_r_1__instr_operands__rs2__18_, calc_stage_r_1__instr_operands__rs2__17_, calc_stage_r_1__instr_operands__rs2__16_, calc_stage_r_1__instr_operands__rs2__15_, calc_stage_r_1__instr_operands__rs2__14_, calc_stage_r_1__instr_operands__rs2__13_, calc_stage_r_1__instr_operands__rs2__12_, calc_stage_r_1__instr_operands__rs2__11_, calc_stage_r_1__instr_operands__rs2__10_, calc_stage_r_1__instr_operands__rs2__9_, calc_stage_r_1__instr_operands__rs2__8_, calc_stage_r_1__instr_operands__rs2__7_, calc_stage_r_1__instr_operands__rs2__6_, calc_stage_r_1__instr_operands__rs2__5_, calc_stage_r_1__instr_operands__rs2__4_, calc_stage_r_1__instr_operands__rs2__3_, calc_stage_r_1__instr_operands__rs2__2_, calc_stage_r_1__instr_operands__rs2__1_, calc_stage_r_1__instr_operands__rs2__0_, calc_stage_r_1__instr_operands__imm__63_, calc_stage_r_1__instr_operands__imm__62_, calc_stage_r_1__instr_operands__imm__61_, calc_stage_r_1__instr_operands__imm__60_, calc_stage_r_1__instr_operands__imm__59_, calc_stage_r_1__instr_operands__imm__58_, calc_stage_r_1__instr_operands__imm__57_, calc_stage_r_1__instr_operands__imm__56_, calc_stage_r_1__instr_operands__imm__55_, calc_stage_r_1__instr_operands__imm__54_, calc_stage_r_1__instr_operands__imm__53_, calc_stage_r_1__instr_operands__imm__52_, calc_stage_r_1__instr_operands__imm__51_, calc_stage_r_1__instr_operands__imm__50_, calc_stage_r_1__instr_operands__imm__49_, calc_stage_r_1__instr_operands__imm__48_, calc_stage_r_1__instr_operands__imm__47_, calc_stage_r_1__instr_operands__imm__46_, calc_stage_r_1__instr_operands__imm__45_, calc_stage_r_1__instr_operands__imm__44_, calc_stage_r_1__instr_operands__imm__43_, calc_stage_r_1__instr_operands__imm__42_, calc_stage_r_1__instr_operands__imm__41_, calc_stage_r_1__instr_operands__imm__40_, calc_stage_r_1__instr_operands__imm__39_, calc_stage_r_1__instr_operands__imm__38_, calc_stage_r_1__instr_operands__imm__37_, calc_stage_r_1__instr_operands__imm__36_, calc_stage_r_1__instr_operands__imm__35_, calc_stage_r_1__instr_operands__imm__34_, calc_stage_r_1__instr_operands__imm__33_, calc_stage_r_1__instr_operands__imm__32_, calc_stage_r_1__instr_operands__imm__31_, calc_stage_r_1__instr_operands__imm__30_, calc_stage_r_1__instr_operands__imm__29_, calc_stage_r_1__instr_operands__imm__28_, calc_stage_r_1__instr_operands__imm__27_, calc_stage_r_1__instr_operands__imm__26_, calc_stage_r_1__instr_operands__imm__25_, calc_stage_r_1__instr_operands__imm__24_, calc_stage_r_1__instr_operands__imm__23_, calc_stage_r_1__instr_operands__imm__22_, calc_stage_r_1__instr_operands__imm__21_, calc_stage_r_1__instr_operands__imm__20_, calc_stage_r_1__instr_operands__imm__19_, calc_stage_r_1__instr_operands__imm__18_, calc_stage_r_1__instr_operands__imm__17_, calc_stage_r_1__instr_operands__imm__16_, calc_stage_r_1__instr_operands__imm__15_, calc_stage_r_1__instr_operands__imm__14_, calc_stage_r_1__instr_operands__imm__13_, calc_stage_r_1__instr_operands__imm__12_, calc_stage_r_1__instr_operands__imm__11_, calc_stage_r_1__instr_operands__imm__10_, calc_stage_r_1__instr_operands__imm__9_, calc_stage_r_1__instr_operands__imm__8_, calc_stage_r_1__instr_operands__imm__7_, calc_stage_r_1__instr_operands__imm__6_, calc_stage_r_1__instr_operands__imm__5_, calc_stage_r_1__instr_operands__imm__4_, calc_stage_r_1__instr_operands__imm__3_, calc_stage_r_1__instr_operands__imm__2_, calc_stage_r_1__instr_operands__imm__1_, calc_stage_r_1__instr_operands__imm__0_, calc_stage_r_1__decode__instr_v_, calc_stage_r_1__decode__fe_nop_v_, calc_stage_r_1__decode__be_nop_v_, calc_stage_r_1__decode__me_nop_v_, calc_stage_r_1__decode__pipe_comp_v_, calc_stage_r_1__decode__pipe_int_v_, calc_stage_r_1__decode__pipe_mul_v_, calc_stage_r_1__decode__pipe_mem_v_, calc_stage_r_1__decode__pipe_fp_v_, calc_stage_r_1__decode__irf_w_v_, calc_stage_r_1__decode__frf_w_v_, calc_stage_r_1__decode__mhartid_r_v_, calc_stage_r_1__decode__dcache_w_v_, calc_stage_r_1__decode__dcache_r_v_, calc_stage_r_1__decode__fp_not_int_v_, calc_stage_r_1__decode__ret_v_, calc_stage_r_1__decode__amo_v_, calc_stage_r_1__decode__jmp_v_, calc_stage_r_1__decode__br_v_, calc_stage_r_1__decode__opw_v_, calc_stage_r_1__decode__fu_op__fu_op__3_, calc_stage_r_1__decode__fu_op__fu_op__2_, calc_stage_r_1__decode__fu_op__fu_op__1_, calc_stage_r_1__decode__fu_op__fu_op__0_, calc_stage_r_1__decode__rs1_addr__4_, calc_stage_r_1__decode__rs1_addr__3_, calc_stage_r_1__decode__rs1_addr__2_, calc_stage_r_1__decode__rs1_addr__1_, calc_stage_r_1__decode__rs1_addr__0_, calc_stage_r_1__decode__rs2_addr__4_, calc_stage_r_1__decode__rs2_addr__3_, calc_stage_r_1__decode__rs2_addr__2_, calc_stage_r_1__decode__rs2_addr__1_, calc_stage_r_1__decode__rs2_addr__0_, calc_status_o[83:79], calc_stage_r_1__decode__src1_sel_, calc_stage_r_1__decode__src2_sel_, calc_stage_r_1__decode__baddr_sel_, calc_stage_r_1__decode__result_sel_, calc_stage_r_0__instr_metadata__itag__7_, calc_stage_r_0__instr_metadata__itag__6_, calc_stage_r_0__instr_metadata__itag__5_, calc_stage_r_0__instr_metadata__itag__4_, calc_stage_r_0__instr_metadata__itag__3_, calc_stage_r_0__instr_metadata__itag__2_, calc_stage_r_0__instr_metadata__itag__1_, calc_stage_r_0__instr_metadata__itag__0_, calc_stage_r_0__instr_metadata__pc__63_, calc_stage_r_0__instr_metadata__pc__62_, calc_stage_r_0__instr_metadata__pc__61_, calc_stage_r_0__instr_metadata__pc__60_, calc_stage_r_0__instr_metadata__pc__59_, calc_stage_r_0__instr_metadata__pc__58_, calc_stage_r_0__instr_metadata__pc__57_, calc_stage_r_0__instr_metadata__pc__56_, calc_stage_r_0__instr_metadata__pc__55_, calc_stage_r_0__instr_metadata__pc__54_, calc_stage_r_0__instr_metadata__pc__53_, calc_stage_r_0__instr_metadata__pc__52_, calc_stage_r_0__instr_metadata__pc__51_, calc_stage_r_0__instr_metadata__pc__50_, calc_stage_r_0__instr_metadata__pc__49_, calc_stage_r_0__instr_metadata__pc__48_, calc_stage_r_0__instr_metadata__pc__47_, calc_stage_r_0__instr_metadata__pc__46_, calc_stage_r_0__instr_metadata__pc__45_, calc_stage_r_0__instr_metadata__pc__44_, calc_stage_r_0__instr_metadata__pc__43_, calc_stage_r_0__instr_metadata__pc__42_, calc_stage_r_0__instr_metadata__pc__41_, calc_stage_r_0__instr_metadata__pc__40_, calc_stage_r_0__instr_metadata__pc__39_, calc_stage_r_0__instr_metadata__pc__38_, calc_stage_r_0__instr_metadata__pc__37_, calc_stage_r_0__instr_metadata__pc__36_, calc_stage_r_0__instr_metadata__pc__35_, calc_stage_r_0__instr_metadata__pc__34_, calc_stage_r_0__instr_metadata__pc__33_, calc_stage_r_0__instr_metadata__pc__32_, calc_stage_r_0__instr_metadata__pc__31_, calc_stage_r_0__instr_metadata__pc__30_, calc_stage_r_0__instr_metadata__pc__29_, calc_stage_r_0__instr_metadata__pc__28_, calc_stage_r_0__instr_metadata__pc__27_, calc_stage_r_0__instr_metadata__pc__26_, calc_stage_r_0__instr_metadata__pc__25_, calc_stage_r_0__instr_metadata__pc__24_, calc_stage_r_0__instr_metadata__pc__23_, calc_stage_r_0__instr_metadata__pc__22_, calc_stage_r_0__instr_metadata__pc__21_, calc_stage_r_0__instr_metadata__pc__20_, calc_stage_r_0__instr_metadata__pc__19_, calc_stage_r_0__instr_metadata__pc__18_, calc_stage_r_0__instr_metadata__pc__17_, calc_stage_r_0__instr_metadata__pc__16_, calc_stage_r_0__instr_metadata__pc__15_, calc_stage_r_0__instr_metadata__pc__14_, calc_stage_r_0__instr_metadata__pc__13_, calc_stage_r_0__instr_metadata__pc__12_, calc_stage_r_0__instr_metadata__pc__11_, calc_stage_r_0__instr_metadata__pc__10_, calc_stage_r_0__instr_metadata__pc__9_, calc_stage_r_0__instr_metadata__pc__8_, calc_stage_r_0__instr_metadata__pc__7_, calc_stage_r_0__instr_metadata__pc__6_, calc_stage_r_0__instr_metadata__pc__5_, calc_stage_r_0__instr_metadata__pc__4_, calc_stage_r_0__instr_metadata__pc__3_, calc_stage_r_0__instr_metadata__pc__2_, calc_stage_r_0__instr_metadata__pc__1_, calc_stage_r_0__instr_metadata__pc__0_, calc_stage_r_0__instr_metadata__fe_exception_not_instr_, calc_stage_r_0__instr_metadata__fe_exception_code__1_, calc_stage_r_0__instr_metadata__fe_exception_code__0_, calc_status_o[157:122], calc_stage_r_0__instr__31_, calc_stage_r_0__instr__30_, calc_stage_r_0__instr__29_, calc_stage_r_0__instr__28_, calc_stage_r_0__instr__27_, calc_stage_r_0__instr__26_, calc_stage_r_0__instr__25_, calc_stage_r_0__instr__24_, calc_stage_r_0__instr__23_, calc_stage_r_0__instr__22_, calc_stage_r_0__instr__21_, calc_stage_r_0__instr__20_, calc_stage_r_0__instr__19_, calc_stage_r_0__instr__18_, calc_stage_r_0__instr__17_, calc_stage_r_0__instr__16_, calc_stage_r_0__instr__15_, calc_stage_r_0__instr__14_, calc_stage_r_0__instr__13_, calc_stage_r_0__instr__12_, calc_stage_r_0__instr__11_, calc_stage_r_0__instr__10_, calc_stage_r_0__instr__9_, calc_stage_r_0__instr__8_, calc_stage_r_0__instr__7_, calc_stage_r_0__instr__6_, calc_stage_r_0__instr__5_, calc_stage_r_0__instr__4_, calc_stage_r_0__instr__3_, calc_stage_r_0__instr__2_, calc_stage_r_0__instr__1_, calc_stage_r_0__instr__0_, calc_stage_r_0__instr_operands__rs1__63_, calc_stage_r_0__instr_operands__rs1__62_, calc_stage_r_0__instr_operands__rs1__61_, calc_stage_r_0__instr_operands__rs1__60_, calc_stage_r_0__instr_operands__rs1__59_, calc_stage_r_0__instr_operands__rs1__58_, calc_stage_r_0__instr_operands__rs1__57_, calc_stage_r_0__instr_operands__rs1__56_, calc_stage_r_0__instr_operands__rs1__55_, calc_stage_r_0__instr_operands__rs1__54_, calc_stage_r_0__instr_operands__rs1__53_, calc_stage_r_0__instr_operands__rs1__52_, calc_stage_r_0__instr_operands__rs1__51_, calc_stage_r_0__instr_operands__rs1__50_, calc_stage_r_0__instr_operands__rs1__49_, calc_stage_r_0__instr_operands__rs1__48_, calc_stage_r_0__instr_operands__rs1__47_, calc_stage_r_0__instr_operands__rs1__46_, calc_stage_r_0__instr_operands__rs1__45_, calc_stage_r_0__instr_operands__rs1__44_, calc_stage_r_0__instr_operands__rs1__43_, calc_stage_r_0__instr_operands__rs1__42_, calc_stage_r_0__instr_operands__rs1__41_, calc_stage_r_0__instr_operands__rs1__40_, calc_stage_r_0__instr_operands__rs1__39_, calc_stage_r_0__instr_operands__rs1__38_, calc_stage_r_0__instr_operands__rs1__37_, calc_stage_r_0__instr_operands__rs1__36_, calc_stage_r_0__instr_operands__rs1__35_, calc_stage_r_0__instr_operands__rs1__34_, calc_stage_r_0__instr_operands__rs1__33_, calc_stage_r_0__instr_operands__rs1__32_, calc_stage_r_0__instr_operands__rs1__31_, calc_stage_r_0__instr_operands__rs1__30_, calc_stage_r_0__instr_operands__rs1__29_, calc_stage_r_0__instr_operands__rs1__28_, calc_stage_r_0__instr_operands__rs1__27_, calc_stage_r_0__instr_operands__rs1__26_, calc_stage_r_0__instr_operands__rs1__25_, calc_stage_r_0__instr_operands__rs1__24_, calc_stage_r_0__instr_operands__rs1__23_, calc_stage_r_0__instr_operands__rs1__22_, calc_stage_r_0__instr_operands__rs1__21_, calc_stage_r_0__instr_operands__rs1__20_, calc_stage_r_0__instr_operands__rs1__19_, calc_stage_r_0__instr_operands__rs1__18_, calc_stage_r_0__instr_operands__rs1__17_, calc_stage_r_0__instr_operands__rs1__16_, calc_stage_r_0__instr_operands__rs1__15_, calc_stage_r_0__instr_operands__rs1__14_, calc_stage_r_0__instr_operands__rs1__13_, calc_stage_r_0__instr_operands__rs1__12_, calc_stage_r_0__instr_operands__rs1__11_, calc_stage_r_0__instr_operands__rs1__10_, calc_stage_r_0__instr_operands__rs1__9_, calc_stage_r_0__instr_operands__rs1__8_, calc_stage_r_0__instr_operands__rs1__7_, calc_stage_r_0__instr_operands__rs1__6_, calc_stage_r_0__instr_operands__rs1__5_, calc_stage_r_0__instr_operands__rs1__4_, calc_stage_r_0__instr_operands__rs1__3_, calc_stage_r_0__instr_operands__rs1__2_, calc_stage_r_0__instr_operands__rs1__1_, calc_stage_r_0__instr_operands__rs1__0_, calc_stage_r_0__instr_operands__rs2__63_, calc_stage_r_0__instr_operands__rs2__62_, calc_stage_r_0__instr_operands__rs2__61_, calc_stage_r_0__instr_operands__rs2__60_, calc_stage_r_0__instr_operands__rs2__59_, calc_stage_r_0__instr_operands__rs2__58_, calc_stage_r_0__instr_operands__rs2__57_, calc_stage_r_0__instr_operands__rs2__56_, calc_stage_r_0__instr_operands__rs2__55_, calc_stage_r_0__instr_operands__rs2__54_, calc_stage_r_0__instr_operands__rs2__53_, calc_stage_r_0__instr_operands__rs2__52_, calc_stage_r_0__instr_operands__rs2__51_, calc_stage_r_0__instr_operands__rs2__50_, calc_stage_r_0__instr_operands__rs2__49_, calc_stage_r_0__instr_operands__rs2__48_, calc_stage_r_0__instr_operands__rs2__47_, calc_stage_r_0__instr_operands__rs2__46_, calc_stage_r_0__instr_operands__rs2__45_, calc_stage_r_0__instr_operands__rs2__44_, calc_stage_r_0__instr_operands__rs2__43_, calc_stage_r_0__instr_operands__rs2__42_, calc_stage_r_0__instr_operands__rs2__41_, calc_stage_r_0__instr_operands__rs2__40_, calc_stage_r_0__instr_operands__rs2__39_, calc_stage_r_0__instr_operands__rs2__38_, calc_stage_r_0__instr_operands__rs2__37_, calc_stage_r_0__instr_operands__rs2__36_, calc_stage_r_0__instr_operands__rs2__35_, calc_stage_r_0__instr_operands__rs2__34_, calc_stage_r_0__instr_operands__rs2__33_, calc_stage_r_0__instr_operands__rs2__32_, calc_stage_r_0__instr_operands__rs2__31_, calc_stage_r_0__instr_operands__rs2__30_, calc_stage_r_0__instr_operands__rs2__29_, calc_stage_r_0__instr_operands__rs2__28_, calc_stage_r_0__instr_operands__rs2__27_, calc_stage_r_0__instr_operands__rs2__26_, calc_stage_r_0__instr_operands__rs2__25_, calc_stage_r_0__instr_operands__rs2__24_, calc_stage_r_0__instr_operands__rs2__23_, calc_stage_r_0__instr_operands__rs2__22_, calc_stage_r_0__instr_operands__rs2__21_, calc_stage_r_0__instr_operands__rs2__20_, calc_stage_r_0__instr_operands__rs2__19_, calc_stage_r_0__instr_operands__rs2__18_, calc_stage_r_0__instr_operands__rs2__17_, calc_stage_r_0__instr_operands__rs2__16_, calc_stage_r_0__instr_operands__rs2__15_, calc_stage_r_0__instr_operands__rs2__14_, calc_stage_r_0__instr_operands__rs2__13_, calc_stage_r_0__instr_operands__rs2__12_, calc_stage_r_0__instr_operands__rs2__11_, calc_stage_r_0__instr_operands__rs2__10_, calc_stage_r_0__instr_operands__rs2__9_, calc_stage_r_0__instr_operands__rs2__8_, calc_stage_r_0__instr_operands__rs2__7_, calc_stage_r_0__instr_operands__rs2__6_, calc_stage_r_0__instr_operands__rs2__5_, calc_stage_r_0__instr_operands__rs2__4_, calc_stage_r_0__instr_operands__rs2__3_, calc_stage_r_0__instr_operands__rs2__2_, calc_stage_r_0__instr_operands__rs2__1_, calc_stage_r_0__instr_operands__rs2__0_, calc_stage_r_0__instr_operands__imm__63_, calc_stage_r_0__instr_operands__imm__62_, calc_stage_r_0__instr_operands__imm__61_, calc_stage_r_0__instr_operands__imm__60_, calc_stage_r_0__instr_operands__imm__59_, calc_stage_r_0__instr_operands__imm__58_, calc_stage_r_0__instr_operands__imm__57_, calc_stage_r_0__instr_operands__imm__56_, calc_stage_r_0__instr_operands__imm__55_, calc_stage_r_0__instr_operands__imm__54_, calc_stage_r_0__instr_operands__imm__53_, calc_stage_r_0__instr_operands__imm__52_, calc_stage_r_0__instr_operands__imm__51_, calc_stage_r_0__instr_operands__imm__50_, calc_stage_r_0__instr_operands__imm__49_, calc_stage_r_0__instr_operands__imm__48_, calc_stage_r_0__instr_operands__imm__47_, calc_stage_r_0__instr_operands__imm__46_, calc_stage_r_0__instr_operands__imm__45_, calc_stage_r_0__instr_operands__imm__44_, calc_stage_r_0__instr_operands__imm__43_, calc_stage_r_0__instr_operands__imm__42_, calc_stage_r_0__instr_operands__imm__41_, calc_stage_r_0__instr_operands__imm__40_, calc_stage_r_0__instr_operands__imm__39_, calc_stage_r_0__instr_operands__imm__38_, calc_stage_r_0__instr_operands__imm__37_, calc_stage_r_0__instr_operands__imm__36_, calc_stage_r_0__instr_operands__imm__35_, calc_stage_r_0__instr_operands__imm__34_, calc_stage_r_0__instr_operands__imm__33_, calc_stage_r_0__instr_operands__imm__32_, calc_stage_r_0__instr_operands__imm__31_, calc_stage_r_0__instr_operands__imm__30_, calc_stage_r_0__instr_operands__imm__29_, calc_stage_r_0__instr_operands__imm__28_, calc_stage_r_0__instr_operands__imm__27_, calc_stage_r_0__instr_operands__imm__26_, calc_stage_r_0__instr_operands__imm__25_, calc_stage_r_0__instr_operands__imm__24_, calc_stage_r_0__instr_operands__imm__23_, calc_stage_r_0__instr_operands__imm__22_, calc_stage_r_0__instr_operands__imm__21_, calc_stage_r_0__instr_operands__imm__20_, calc_stage_r_0__instr_operands__imm__19_, calc_stage_r_0__instr_operands__imm__18_, calc_stage_r_0__instr_operands__imm__17_, calc_stage_r_0__instr_operands__imm__16_, calc_stage_r_0__instr_operands__imm__15_, calc_stage_r_0__instr_operands__imm__14_, calc_stage_r_0__instr_operands__imm__13_, calc_stage_r_0__instr_operands__imm__12_, calc_stage_r_0__instr_operands__imm__11_, calc_stage_r_0__instr_operands__imm__10_, calc_stage_r_0__instr_operands__imm__9_, calc_stage_r_0__instr_operands__imm__8_, calc_stage_r_0__instr_operands__imm__7_, calc_stage_r_0__instr_operands__imm__6_, calc_stage_r_0__instr_operands__imm__5_, calc_stage_r_0__instr_operands__imm__4_, calc_stage_r_0__instr_operands__imm__3_, calc_stage_r_0__instr_operands__imm__2_, calc_stage_r_0__instr_operands__imm__1_, calc_stage_r_0__instr_operands__imm__0_, calc_stage_r_0__decode__instr_v_, calc_stage_r_0__decode__fe_nop_v_, calc_stage_r_0__decode__be_nop_v_, calc_stage_r_0__decode__me_nop_v_, calc_stage_r_0__decode__pipe_comp_v_, calc_stage_r_0__decode__pipe_int_v_, calc_stage_r_0__decode__pipe_mul_v_, calc_stage_r_0__decode__pipe_mem_v_, calc_stage_r_0__decode__pipe_fp_v_, calc_stage_r_0__decode__irf_w_v_, calc_stage_r_0__decode__frf_w_v_, calc_stage_r_0__decode__mhartid_r_v_, calc_stage_r_0__decode__dcache_w_v_, calc_stage_r_0__decode__dcache_r_v_, calc_stage_r_0__decode__fp_not_int_v_, calc_stage_r_0__decode__ret_v_, calc_stage_r_0__decode__amo_v_, calc_stage_r_0__decode__jmp_v_, calc_stage_r_0__decode__br_v_, calc_stage_r_0__decode__opw_v_, calc_stage_r_0__decode__fu_op__fu_op__3_, calc_stage_r_0__decode__fu_op__fu_op__2_, calc_stage_r_0__decode__fu_op__fu_op__1_, calc_stage_r_0__decode__fu_op__fu_op__0_, calc_stage_r_0__decode__rs1_addr__4_, calc_stage_r_0__decode__rs1_addr__3_, calc_stage_r_0__decode__rs1_addr__2_, calc_stage_r_0__decode__rs1_addr__1_, calc_stage_r_0__decode__rs1_addr__0_, calc_stage_r_0__decode__rs2_addr__4_, calc_stage_r_0__decode__rs2_addr__3_, calc_stage_r_0__decode__rs2_addr__2_, calc_stage_r_0__decode__rs2_addr__1_, calc_stage_r_0__decode__rs2_addr__0_, calc_status_o[73:69], calc_stage_r_0__decode__src1_sel_, calc_stage_r_0__decode__src2_sel_, calc_stage_r_0__decode__baddr_sel_, calc_stage_r_0__decode__result_sel_, dispatch_pkt_instr_metadata__itag__7_, dispatch_pkt_instr_metadata__itag__6_, dispatch_pkt_instr_metadata__itag__5_, dispatch_pkt_instr_metadata__itag__4_, dispatch_pkt_instr_metadata__itag__3_, dispatch_pkt_instr_metadata__itag__2_, dispatch_pkt_instr_metadata__itag__1_, dispatch_pkt_instr_metadata__itag__0_, calc_status_o[300:237], dispatch_pkt_instr_metadata__fe_exception_not_instr_, dispatch_pkt_instr_metadata__fe_exception_code__1_, dispatch_pkt_instr_metadata__fe_exception_code__0_, dispatch_pkt_instr_metadata__branch_metadata_fwd__35_, dispatch_pkt_instr_metadata__branch_metadata_fwd__34_, dispatch_pkt_instr_metadata__branch_metadata_fwd__33_, dispatch_pkt_instr_metadata__branch_metadata_fwd__32_, dispatch_pkt_instr_metadata__branch_metadata_fwd__31_, dispatch_pkt_instr_metadata__branch_metadata_fwd__30_, dispatch_pkt_instr_metadata__branch_metadata_fwd__29_, dispatch_pkt_instr_metadata__branch_metadata_fwd__28_, dispatch_pkt_instr_metadata__branch_metadata_fwd__27_, dispatch_pkt_instr_metadata__branch_metadata_fwd__26_, dispatch_pkt_instr_metadata__branch_metadata_fwd__25_, dispatch_pkt_instr_metadata__branch_metadata_fwd__24_, dispatch_pkt_instr_metadata__branch_metadata_fwd__23_, dispatch_pkt_instr_metadata__branch_metadata_fwd__22_, dispatch_pkt_instr_metadata__branch_metadata_fwd__21_, dispatch_pkt_instr_metadata__branch_metadata_fwd__20_, dispatch_pkt_instr_metadata__branch_metadata_fwd__19_, dispatch_pkt_instr_metadata__branch_metadata_fwd__18_, dispatch_pkt_instr_metadata__branch_metadata_fwd__17_, dispatch_pkt_instr_metadata__branch_metadata_fwd__16_, dispatch_pkt_instr_metadata__branch_metadata_fwd__15_, dispatch_pkt_instr_metadata__branch_metadata_fwd__14_, dispatch_pkt_instr_metadata__branch_metadata_fwd__13_, dispatch_pkt_instr_metadata__branch_metadata_fwd__12_, dispatch_pkt_instr_metadata__branch_metadata_fwd__11_, dispatch_pkt_instr_metadata__branch_metadata_fwd__10_, dispatch_pkt_instr_metadata__branch_metadata_fwd__9_, dispatch_pkt_instr_metadata__branch_metadata_fwd__8_, dispatch_pkt_instr_metadata__branch_metadata_fwd__7_, dispatch_pkt_instr_metadata__branch_metadata_fwd__6_, dispatch_pkt_instr_metadata__branch_metadata_fwd__5_, dispatch_pkt_instr_metadata__branch_metadata_fwd__4_, dispatch_pkt_instr_metadata__branch_metadata_fwd__3_, dispatch_pkt_instr_metadata__branch_metadata_fwd__2_, dispatch_pkt_instr_metadata__branch_metadata_fwd__1_, dispatch_pkt_instr_metadata__branch_metadata_fwd__0_, issue_pkt_r_instr__31_, issue_pkt_r_instr__30_, issue_pkt_r_instr__29_, issue_pkt_r_instr__28_, issue_pkt_r_instr__27_, issue_pkt_r_instr__26_, issue_pkt_r_instr__25_, issue_pkt_r_instr__24_, issue_pkt_r_instr__23_, issue_pkt_r_instr__22_, issue_pkt_r_instr__21_, issue_pkt_r_instr__20_, issue_pkt_r_instr__19_, issue_pkt_r_instr__18_, issue_pkt_r_instr__17_, issue_pkt_r_instr__16_, issue_pkt_r_instr__15_, issue_pkt_r_instr__14_, issue_pkt_r_instr__13_, issue_pkt_r_instr__12_, issue_pkt_r_instr__11_, issue_pkt_r_instr__10_, issue_pkt_r_instr__9_, issue_pkt_r_instr__8_, issue_pkt_r_instr__7_, issue_pkt_r_instr__6_, issue_pkt_r_instr__5_, issue_pkt_r_instr__4_, issue_pkt_r_instr__3_, issue_pkt_r_instr__2_, issue_pkt_r_instr__1_, issue_pkt_r_instr__0_, dispatch_pkt_instr_operands__rs1__63_, dispatch_pkt_instr_operands__rs1__62_, dispatch_pkt_instr_operands__rs1__61_, dispatch_pkt_instr_operands__rs1__60_, dispatch_pkt_instr_operands__rs1__59_, dispatch_pkt_instr_operands__rs1__58_, dispatch_pkt_instr_operands__rs1__57_, dispatch_pkt_instr_operands__rs1__56_, dispatch_pkt_instr_operands__rs1__55_, dispatch_pkt_instr_operands__rs1__54_, dispatch_pkt_instr_operands__rs1__53_, dispatch_pkt_instr_operands__rs1__52_, dispatch_pkt_instr_operands__rs1__51_, dispatch_pkt_instr_operands__rs1__50_, dispatch_pkt_instr_operands__rs1__49_, dispatch_pkt_instr_operands__rs1__48_, dispatch_pkt_instr_operands__rs1__47_, dispatch_pkt_instr_operands__rs1__46_, dispatch_pkt_instr_operands__rs1__45_, dispatch_pkt_instr_operands__rs1__44_, dispatch_pkt_instr_operands__rs1__43_, dispatch_pkt_instr_operands__rs1__42_, dispatch_pkt_instr_operands__rs1__41_, dispatch_pkt_instr_operands__rs1__40_, dispatch_pkt_instr_operands__rs1__39_, dispatch_pkt_instr_operands__rs1__38_, dispatch_pkt_instr_operands__rs1__37_, dispatch_pkt_instr_operands__rs1__36_, dispatch_pkt_instr_operands__rs1__35_, dispatch_pkt_instr_operands__rs1__34_, dispatch_pkt_instr_operands__rs1__33_, dispatch_pkt_instr_operands__rs1__32_, dispatch_pkt_instr_operands__rs1__31_, dispatch_pkt_instr_operands__rs1__30_, dispatch_pkt_instr_operands__rs1__29_, dispatch_pkt_instr_operands__rs1__28_, dispatch_pkt_instr_operands__rs1__27_, dispatch_pkt_instr_operands__rs1__26_, dispatch_pkt_instr_operands__rs1__25_, dispatch_pkt_instr_operands__rs1__24_, dispatch_pkt_instr_operands__rs1__23_, dispatch_pkt_instr_operands__rs1__22_, dispatch_pkt_instr_operands__rs1__21_, dispatch_pkt_instr_operands__rs1__20_, dispatch_pkt_instr_operands__rs1__19_, dispatch_pkt_instr_operands__rs1__18_, dispatch_pkt_instr_operands__rs1__17_, dispatch_pkt_instr_operands__rs1__16_, dispatch_pkt_instr_operands__rs1__15_, dispatch_pkt_instr_operands__rs1__14_, dispatch_pkt_instr_operands__rs1__13_, dispatch_pkt_instr_operands__rs1__12_, dispatch_pkt_instr_operands__rs1__11_, dispatch_pkt_instr_operands__rs1__10_, dispatch_pkt_instr_operands__rs1__9_, dispatch_pkt_instr_operands__rs1__8_, dispatch_pkt_instr_operands__rs1__7_, dispatch_pkt_instr_operands__rs1__6_, dispatch_pkt_instr_operands__rs1__5_, dispatch_pkt_instr_operands__rs1__4_, dispatch_pkt_instr_operands__rs1__3_, dispatch_pkt_instr_operands__rs1__2_, dispatch_pkt_instr_operands__rs1__1_, dispatch_pkt_instr_operands__rs1__0_, dispatch_pkt_instr_operands__rs2__63_, dispatch_pkt_instr_operands__rs2__62_, dispatch_pkt_instr_operands__rs2__61_, dispatch_pkt_instr_operands__rs2__60_, dispatch_pkt_instr_operands__rs2__59_, dispatch_pkt_instr_operands__rs2__58_, dispatch_pkt_instr_operands__rs2__57_, dispatch_pkt_instr_operands__rs2__56_, dispatch_pkt_instr_operands__rs2__55_, dispatch_pkt_instr_operands__rs2__54_, dispatch_pkt_instr_operands__rs2__53_, dispatch_pkt_instr_operands__rs2__52_, dispatch_pkt_instr_operands__rs2__51_, dispatch_pkt_instr_operands__rs2__50_, dispatch_pkt_instr_operands__rs2__49_, dispatch_pkt_instr_operands__rs2__48_, dispatch_pkt_instr_operands__rs2__47_, dispatch_pkt_instr_operands__rs2__46_, dispatch_pkt_instr_operands__rs2__45_, dispatch_pkt_instr_operands__rs2__44_, dispatch_pkt_instr_operands__rs2__43_, dispatch_pkt_instr_operands__rs2__42_, dispatch_pkt_instr_operands__rs2__41_, dispatch_pkt_instr_operands__rs2__40_, dispatch_pkt_instr_operands__rs2__39_, dispatch_pkt_instr_operands__rs2__38_, dispatch_pkt_instr_operands__rs2__37_, dispatch_pkt_instr_operands__rs2__36_, dispatch_pkt_instr_operands__rs2__35_, dispatch_pkt_instr_operands__rs2__34_, dispatch_pkt_instr_operands__rs2__33_, dispatch_pkt_instr_operands__rs2__32_, dispatch_pkt_instr_operands__rs2__31_, dispatch_pkt_instr_operands__rs2__30_, dispatch_pkt_instr_operands__rs2__29_, dispatch_pkt_instr_operands__rs2__28_, dispatch_pkt_instr_operands__rs2__27_, dispatch_pkt_instr_operands__rs2__26_, dispatch_pkt_instr_operands__rs2__25_, dispatch_pkt_instr_operands__rs2__24_, dispatch_pkt_instr_operands__rs2__23_, dispatch_pkt_instr_operands__rs2__22_, dispatch_pkt_instr_operands__rs2__21_, dispatch_pkt_instr_operands__rs2__20_, dispatch_pkt_instr_operands__rs2__19_, dispatch_pkt_instr_operands__rs2__18_, dispatch_pkt_instr_operands__rs2__17_, dispatch_pkt_instr_operands__rs2__16_, dispatch_pkt_instr_operands__rs2__15_, dispatch_pkt_instr_operands__rs2__14_, dispatch_pkt_instr_operands__rs2__13_, dispatch_pkt_instr_operands__rs2__12_, dispatch_pkt_instr_operands__rs2__11_, dispatch_pkt_instr_operands__rs2__10_, dispatch_pkt_instr_operands__rs2__9_, dispatch_pkt_instr_operands__rs2__8_, dispatch_pkt_instr_operands__rs2__7_, dispatch_pkt_instr_operands__rs2__6_, dispatch_pkt_instr_operands__rs2__5_, dispatch_pkt_instr_operands__rs2__4_, dispatch_pkt_instr_operands__rs2__3_, dispatch_pkt_instr_operands__rs2__2_, dispatch_pkt_instr_operands__rs2__1_, dispatch_pkt_instr_operands__rs2__0_, dispatch_pkt_instr_operands__imm__63_, dispatch_pkt_instr_operands__imm__62_, dispatch_pkt_instr_operands__imm__61_, dispatch_pkt_instr_operands__imm__60_, dispatch_pkt_instr_operands__imm__59_, dispatch_pkt_instr_operands__imm__58_, dispatch_pkt_instr_operands__imm__57_, dispatch_pkt_instr_operands__imm__56_, dispatch_pkt_instr_operands__imm__55_, dispatch_pkt_instr_operands__imm__54_, dispatch_pkt_instr_operands__imm__53_, dispatch_pkt_instr_operands__imm__52_, dispatch_pkt_instr_operands__imm__51_, dispatch_pkt_instr_operands__imm__50_, dispatch_pkt_instr_operands__imm__49_, dispatch_pkt_instr_operands__imm__48_, dispatch_pkt_instr_operands__imm__47_, dispatch_pkt_instr_operands__imm__46_, dispatch_pkt_instr_operands__imm__45_, dispatch_pkt_instr_operands__imm__44_, dispatch_pkt_instr_operands__imm__43_, dispatch_pkt_instr_operands__imm__42_, dispatch_pkt_instr_operands__imm__41_, dispatch_pkt_instr_operands__imm__40_, dispatch_pkt_instr_operands__imm__39_, dispatch_pkt_instr_operands__imm__38_, dispatch_pkt_instr_operands__imm__37_, dispatch_pkt_instr_operands__imm__36_, dispatch_pkt_instr_operands__imm__35_, dispatch_pkt_instr_operands__imm__34_, dispatch_pkt_instr_operands__imm__33_, dispatch_pkt_instr_operands__imm__32_, dispatch_pkt_instr_operands__imm__31_, dispatch_pkt_instr_operands__imm__30_, dispatch_pkt_instr_operands__imm__29_, dispatch_pkt_instr_operands__imm__28_, dispatch_pkt_instr_operands__imm__27_, dispatch_pkt_instr_operands__imm__26_, dispatch_pkt_instr_operands__imm__25_, dispatch_pkt_instr_operands__imm__24_, dispatch_pkt_instr_operands__imm__23_, dispatch_pkt_instr_operands__imm__22_, dispatch_pkt_instr_operands__imm__21_, dispatch_pkt_instr_operands__imm__20_, dispatch_pkt_instr_operands__imm__19_, dispatch_pkt_instr_operands__imm__18_, dispatch_pkt_instr_operands__imm__17_, dispatch_pkt_instr_operands__imm__16_, dispatch_pkt_instr_operands__imm__15_, dispatch_pkt_instr_operands__imm__14_, dispatch_pkt_instr_operands__imm__13_, dispatch_pkt_instr_operands__imm__12_, dispatch_pkt_instr_operands__imm__11_, dispatch_pkt_instr_operands__imm__10_, dispatch_pkt_instr_operands__imm__9_, dispatch_pkt_instr_operands__imm__8_, dispatch_pkt_instr_operands__imm__7_, dispatch_pkt_instr_operands__imm__6_, dispatch_pkt_instr_operands__imm__5_, dispatch_pkt_instr_operands__imm__4_, dispatch_pkt_instr_operands__imm__3_, dispatch_pkt_instr_operands__imm__2_, dispatch_pkt_instr_operands__imm__1_, dispatch_pkt_instr_operands__imm__0_, dispatch_pkt_decode__instr_v_, dispatch_pkt_decode__fe_nop_v_, dispatch_pkt_decode__be_nop_v_, dispatch_pkt_decode__me_nop_v_, dispatch_pkt_decode__pipe_comp_v_, dispatch_pkt_decode__pipe_int_v_, dispatch_pkt_decode__pipe_mul_v_, dispatch_pkt_decode__pipe_mem_v_, dispatch_pkt_decode__pipe_fp_v_, dispatch_pkt_decode__irf_w_v_, dispatch_pkt_decode__frf_w_v_, dispatch_pkt_decode__mhartid_r_v_, dispatch_pkt_decode__dcache_w_v_, dispatch_pkt_decode__dcache_r_v_, decoded_fp_not_int_v_, dispatch_pkt_decode__ret_v_, dispatch_pkt_decode__amo_v_, dispatch_pkt_decode__jmp_v_, dispatch_pkt_decode__br_v_, dispatch_pkt_decode__opw_v_, decoded_fu_op_o, decoded_rs1_addr__4_, decoded_rs1_addr__3_, decoded_rs1_addr__2_, decoded_rs1_addr__1_, decoded_rs1_addr__0_, decoded_rs2_addr__4_, decoded_rs2_addr__3_, decoded_rs2_addr__2_, decoded_rs2_addr__1_, decoded_rs2_addr__0_, dispatch_pkt_decode__rd_addr__4_, dispatch_pkt_decode__rd_addr__3_, dispatch_pkt_decode__rd_addr__2_, dispatch_pkt_decode__rd_addr__1_, dispatch_pkt_decode__rd_addr__0_, dispatch_pkt_decode__src1_sel_, dispatch_pkt_decode__src2_sel_, dispatch_pkt_decode__baddr_sel_, dispatch_pkt_decode__result_sel_ }),
    .data_o({ cmt_trace_stage_reg_o[377:9], calc_status_o[113:109], cmt_trace_stage_reg_o[3:0], calc_stage_r_3__instr_metadata__itag__7_, calc_stage_r_3__instr_metadata__itag__6_, calc_stage_r_3__instr_metadata__itag__5_, calc_stage_r_3__instr_metadata__itag__4_, calc_stage_r_3__instr_metadata__itag__3_, calc_stage_r_3__instr_metadata__itag__2_, calc_stage_r_3__instr_metadata__itag__1_, calc_stage_r_3__instr_metadata__itag__0_, calc_stage_r_3__instr_metadata__pc__63_, calc_stage_r_3__instr_metadata__pc__62_, calc_stage_r_3__instr_metadata__pc__61_, calc_stage_r_3__instr_metadata__pc__60_, calc_stage_r_3__instr_metadata__pc__59_, calc_stage_r_3__instr_metadata__pc__58_, calc_stage_r_3__instr_metadata__pc__57_, calc_stage_r_3__instr_metadata__pc__56_, calc_stage_r_3__instr_metadata__pc__55_, calc_stage_r_3__instr_metadata__pc__54_, calc_stage_r_3__instr_metadata__pc__53_, calc_stage_r_3__instr_metadata__pc__52_, calc_stage_r_3__instr_metadata__pc__51_, calc_stage_r_3__instr_metadata__pc__50_, calc_stage_r_3__instr_metadata__pc__49_, calc_stage_r_3__instr_metadata__pc__48_, calc_stage_r_3__instr_metadata__pc__47_, calc_stage_r_3__instr_metadata__pc__46_, calc_stage_r_3__instr_metadata__pc__45_, calc_stage_r_3__instr_metadata__pc__44_, calc_stage_r_3__instr_metadata__pc__43_, calc_stage_r_3__instr_metadata__pc__42_, calc_stage_r_3__instr_metadata__pc__41_, calc_stage_r_3__instr_metadata__pc__40_, calc_stage_r_3__instr_metadata__pc__39_, calc_stage_r_3__instr_metadata__pc__38_, calc_stage_r_3__instr_metadata__pc__37_, calc_stage_r_3__instr_metadata__pc__36_, calc_stage_r_3__instr_metadata__pc__35_, calc_stage_r_3__instr_metadata__pc__34_, calc_stage_r_3__instr_metadata__pc__33_, calc_stage_r_3__instr_metadata__pc__32_, calc_stage_r_3__instr_metadata__pc__31_, calc_stage_r_3__instr_metadata__pc__30_, calc_stage_r_3__instr_metadata__pc__29_, calc_stage_r_3__instr_metadata__pc__28_, calc_stage_r_3__instr_metadata__pc__27_, calc_stage_r_3__instr_metadata__pc__26_, calc_stage_r_3__instr_metadata__pc__25_, calc_stage_r_3__instr_metadata__pc__24_, calc_stage_r_3__instr_metadata__pc__23_, calc_stage_r_3__instr_metadata__pc__22_, calc_stage_r_3__instr_metadata__pc__21_, calc_stage_r_3__instr_metadata__pc__20_, calc_stage_r_3__instr_metadata__pc__19_, calc_stage_r_3__instr_metadata__pc__18_, calc_stage_r_3__instr_metadata__pc__17_, calc_stage_r_3__instr_metadata__pc__16_, calc_stage_r_3__instr_metadata__pc__15_, calc_stage_r_3__instr_metadata__pc__14_, calc_stage_r_3__instr_metadata__pc__13_, calc_stage_r_3__instr_metadata__pc__12_, calc_stage_r_3__instr_metadata__pc__11_, calc_stage_r_3__instr_metadata__pc__10_, calc_stage_r_3__instr_metadata__pc__9_, calc_stage_r_3__instr_metadata__pc__8_, calc_stage_r_3__instr_metadata__pc__7_, calc_stage_r_3__instr_metadata__pc__6_, calc_stage_r_3__instr_metadata__pc__5_, calc_stage_r_3__instr_metadata__pc__4_, calc_stage_r_3__instr_metadata__pc__3_, calc_stage_r_3__instr_metadata__pc__2_, calc_stage_r_3__instr_metadata__pc__1_, calc_stage_r_3__instr_metadata__pc__0_, calc_stage_r_3__instr_metadata__fe_exception_not_instr_, calc_stage_r_3__instr_metadata__fe_exception_code__1_, calc_stage_r_3__instr_metadata__fe_exception_code__0_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__35_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__34_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__33_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__32_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__31_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__30_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__29_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__28_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__27_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__26_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__25_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__24_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__23_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__22_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__21_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__20_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__19_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__18_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__17_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__16_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__15_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__14_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__13_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__12_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__11_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__10_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__9_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__8_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__7_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__6_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__5_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__4_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__3_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__2_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__1_, calc_stage_r_3__instr_metadata__branch_metadata_fwd__0_, calc_stage_r_3__instr__31_, calc_stage_r_3__instr__30_, calc_stage_r_3__instr__29_, calc_stage_r_3__instr__28_, calc_stage_r_3__instr__27_, calc_stage_r_3__instr__26_, calc_stage_r_3__instr__25_, calc_stage_r_3__instr__24_, calc_stage_r_3__instr__23_, calc_stage_r_3__instr__22_, calc_stage_r_3__instr__21_, calc_stage_r_3__instr__20_, calc_stage_r_3__instr__19_, calc_stage_r_3__instr__18_, calc_stage_r_3__instr__17_, calc_stage_r_3__instr__16_, calc_stage_r_3__instr__15_, calc_stage_r_3__instr__14_, calc_stage_r_3__instr__13_, calc_stage_r_3__instr__12_, calc_stage_r_3__instr__11_, calc_stage_r_3__instr__10_, calc_stage_r_3__instr__9_, calc_stage_r_3__instr__8_, calc_stage_r_3__instr__7_, calc_stage_r_3__instr__6_, calc_stage_r_3__instr__5_, calc_stage_r_3__instr__4_, calc_stage_r_3__instr__3_, calc_stage_r_3__instr__2_, calc_stage_r_3__instr__1_, calc_stage_r_3__instr__0_, calc_stage_r_3__instr_operands__rs1__63_, calc_stage_r_3__instr_operands__rs1__62_, calc_stage_r_3__instr_operands__rs1__61_, calc_stage_r_3__instr_operands__rs1__60_, calc_stage_r_3__instr_operands__rs1__59_, calc_stage_r_3__instr_operands__rs1__58_, calc_stage_r_3__instr_operands__rs1__57_, calc_stage_r_3__instr_operands__rs1__56_, calc_stage_r_3__instr_operands__rs1__55_, calc_stage_r_3__instr_operands__rs1__54_, calc_stage_r_3__instr_operands__rs1__53_, calc_stage_r_3__instr_operands__rs1__52_, calc_stage_r_3__instr_operands__rs1__51_, calc_stage_r_3__instr_operands__rs1__50_, calc_stage_r_3__instr_operands__rs1__49_, calc_stage_r_3__instr_operands__rs1__48_, calc_stage_r_3__instr_operands__rs1__47_, calc_stage_r_3__instr_operands__rs1__46_, calc_stage_r_3__instr_operands__rs1__45_, calc_stage_r_3__instr_operands__rs1__44_, calc_stage_r_3__instr_operands__rs1__43_, calc_stage_r_3__instr_operands__rs1__42_, calc_stage_r_3__instr_operands__rs1__41_, calc_stage_r_3__instr_operands__rs1__40_, calc_stage_r_3__instr_operands__rs1__39_, calc_stage_r_3__instr_operands__rs1__38_, calc_stage_r_3__instr_operands__rs1__37_, calc_stage_r_3__instr_operands__rs1__36_, calc_stage_r_3__instr_operands__rs1__35_, calc_stage_r_3__instr_operands__rs1__34_, calc_stage_r_3__instr_operands__rs1__33_, calc_stage_r_3__instr_operands__rs1__32_, calc_stage_r_3__instr_operands__rs1__31_, calc_stage_r_3__instr_operands__rs1__30_, calc_stage_r_3__instr_operands__rs1__29_, calc_stage_r_3__instr_operands__rs1__28_, calc_stage_r_3__instr_operands__rs1__27_, calc_stage_r_3__instr_operands__rs1__26_, calc_stage_r_3__instr_operands__rs1__25_, calc_stage_r_3__instr_operands__rs1__24_, calc_stage_r_3__instr_operands__rs1__23_, calc_stage_r_3__instr_operands__rs1__22_, calc_stage_r_3__instr_operands__rs1__21_, calc_stage_r_3__instr_operands__rs1__20_, calc_stage_r_3__instr_operands__rs1__19_, calc_stage_r_3__instr_operands__rs1__18_, calc_stage_r_3__instr_operands__rs1__17_, calc_stage_r_3__instr_operands__rs1__16_, calc_stage_r_3__instr_operands__rs1__15_, calc_stage_r_3__instr_operands__rs1__14_, calc_stage_r_3__instr_operands__rs1__13_, calc_stage_r_3__instr_operands__rs1__12_, calc_stage_r_3__instr_operands__rs1__11_, calc_stage_r_3__instr_operands__rs1__10_, calc_stage_r_3__instr_operands__rs1__9_, calc_stage_r_3__instr_operands__rs1__8_, calc_stage_r_3__instr_operands__rs1__7_, calc_stage_r_3__instr_operands__rs1__6_, calc_stage_r_3__instr_operands__rs1__5_, calc_stage_r_3__instr_operands__rs1__4_, calc_stage_r_3__instr_operands__rs1__3_, calc_stage_r_3__instr_operands__rs1__2_, calc_stage_r_3__instr_operands__rs1__1_, calc_stage_r_3__instr_operands__rs1__0_, calc_stage_r_3__instr_operands__rs2__63_, calc_stage_r_3__instr_operands__rs2__62_, calc_stage_r_3__instr_operands__rs2__61_, calc_stage_r_3__instr_operands__rs2__60_, calc_stage_r_3__instr_operands__rs2__59_, calc_stage_r_3__instr_operands__rs2__58_, calc_stage_r_3__instr_operands__rs2__57_, calc_stage_r_3__instr_operands__rs2__56_, calc_stage_r_3__instr_operands__rs2__55_, calc_stage_r_3__instr_operands__rs2__54_, calc_stage_r_3__instr_operands__rs2__53_, calc_stage_r_3__instr_operands__rs2__52_, calc_stage_r_3__instr_operands__rs2__51_, calc_stage_r_3__instr_operands__rs2__50_, calc_stage_r_3__instr_operands__rs2__49_, calc_stage_r_3__instr_operands__rs2__48_, calc_stage_r_3__instr_operands__rs2__47_, calc_stage_r_3__instr_operands__rs2__46_, calc_stage_r_3__instr_operands__rs2__45_, calc_stage_r_3__instr_operands__rs2__44_, calc_stage_r_3__instr_operands__rs2__43_, calc_stage_r_3__instr_operands__rs2__42_, calc_stage_r_3__instr_operands__rs2__41_, calc_stage_r_3__instr_operands__rs2__40_, calc_stage_r_3__instr_operands__rs2__39_, calc_stage_r_3__instr_operands__rs2__38_, calc_stage_r_3__instr_operands__rs2__37_, calc_stage_r_3__instr_operands__rs2__36_, calc_stage_r_3__instr_operands__rs2__35_, calc_stage_r_3__instr_operands__rs2__34_, calc_stage_r_3__instr_operands__rs2__33_, calc_stage_r_3__instr_operands__rs2__32_, calc_stage_r_3__instr_operands__rs2__31_, calc_stage_r_3__instr_operands__rs2__30_, calc_stage_r_3__instr_operands__rs2__29_, calc_stage_r_3__instr_operands__rs2__28_, calc_stage_r_3__instr_operands__rs2__27_, calc_stage_r_3__instr_operands__rs2__26_, calc_stage_r_3__instr_operands__rs2__25_, calc_stage_r_3__instr_operands__rs2__24_, calc_stage_r_3__instr_operands__rs2__23_, calc_stage_r_3__instr_operands__rs2__22_, calc_stage_r_3__instr_operands__rs2__21_, calc_stage_r_3__instr_operands__rs2__20_, calc_stage_r_3__instr_operands__rs2__19_, calc_stage_r_3__instr_operands__rs2__18_, calc_stage_r_3__instr_operands__rs2__17_, calc_stage_r_3__instr_operands__rs2__16_, calc_stage_r_3__instr_operands__rs2__15_, calc_stage_r_3__instr_operands__rs2__14_, calc_stage_r_3__instr_operands__rs2__13_, calc_stage_r_3__instr_operands__rs2__12_, calc_stage_r_3__instr_operands__rs2__11_, calc_stage_r_3__instr_operands__rs2__10_, calc_stage_r_3__instr_operands__rs2__9_, calc_stage_r_3__instr_operands__rs2__8_, calc_stage_r_3__instr_operands__rs2__7_, calc_stage_r_3__instr_operands__rs2__6_, calc_stage_r_3__instr_operands__rs2__5_, calc_stage_r_3__instr_operands__rs2__4_, calc_stage_r_3__instr_operands__rs2__3_, calc_stage_r_3__instr_operands__rs2__2_, calc_stage_r_3__instr_operands__rs2__1_, calc_stage_r_3__instr_operands__rs2__0_, calc_stage_r_3__instr_operands__imm__63_, calc_stage_r_3__instr_operands__imm__62_, calc_stage_r_3__instr_operands__imm__61_, calc_stage_r_3__instr_operands__imm__60_, calc_stage_r_3__instr_operands__imm__59_, calc_stage_r_3__instr_operands__imm__58_, calc_stage_r_3__instr_operands__imm__57_, calc_stage_r_3__instr_operands__imm__56_, calc_stage_r_3__instr_operands__imm__55_, calc_stage_r_3__instr_operands__imm__54_, calc_stage_r_3__instr_operands__imm__53_, calc_stage_r_3__instr_operands__imm__52_, calc_stage_r_3__instr_operands__imm__51_, calc_stage_r_3__instr_operands__imm__50_, calc_stage_r_3__instr_operands__imm__49_, calc_stage_r_3__instr_operands__imm__48_, calc_stage_r_3__instr_operands__imm__47_, calc_stage_r_3__instr_operands__imm__46_, calc_stage_r_3__instr_operands__imm__45_, calc_stage_r_3__instr_operands__imm__44_, calc_stage_r_3__instr_operands__imm__43_, calc_stage_r_3__instr_operands__imm__42_, calc_stage_r_3__instr_operands__imm__41_, calc_stage_r_3__instr_operands__imm__40_, calc_stage_r_3__instr_operands__imm__39_, calc_stage_r_3__instr_operands__imm__38_, calc_stage_r_3__instr_operands__imm__37_, calc_stage_r_3__instr_operands__imm__36_, calc_stage_r_3__instr_operands__imm__35_, calc_stage_r_3__instr_operands__imm__34_, calc_stage_r_3__instr_operands__imm__33_, calc_stage_r_3__instr_operands__imm__32_, calc_stage_r_3__instr_operands__imm__31_, calc_stage_r_3__instr_operands__imm__30_, calc_stage_r_3__instr_operands__imm__29_, calc_stage_r_3__instr_operands__imm__28_, calc_stage_r_3__instr_operands__imm__27_, calc_stage_r_3__instr_operands__imm__26_, calc_stage_r_3__instr_operands__imm__25_, calc_stage_r_3__instr_operands__imm__24_, calc_stage_r_3__instr_operands__imm__23_, calc_stage_r_3__instr_operands__imm__22_, calc_stage_r_3__instr_operands__imm__21_, calc_stage_r_3__instr_operands__imm__20_, calc_stage_r_3__instr_operands__imm__19_, calc_stage_r_3__instr_operands__imm__18_, calc_stage_r_3__instr_operands__imm__17_, calc_stage_r_3__instr_operands__imm__16_, calc_stage_r_3__instr_operands__imm__15_, calc_stage_r_3__instr_operands__imm__14_, calc_stage_r_3__instr_operands__imm__13_, calc_stage_r_3__instr_operands__imm__12_, calc_stage_r_3__instr_operands__imm__11_, calc_stage_r_3__instr_operands__imm__10_, calc_stage_r_3__instr_operands__imm__9_, calc_stage_r_3__instr_operands__imm__8_, calc_stage_r_3__instr_operands__imm__7_, calc_stage_r_3__instr_operands__imm__6_, calc_stage_r_3__instr_operands__imm__5_, calc_stage_r_3__instr_operands__imm__4_, calc_stage_r_3__instr_operands__imm__3_, calc_stage_r_3__instr_operands__imm__2_, calc_stage_r_3__instr_operands__imm__1_, calc_stage_r_3__instr_operands__imm__0_, calc_stage_r_3__decode__instr_v_, calc_stage_r_3__decode__fe_nop_v_, calc_stage_r_3__decode__be_nop_v_, calc_stage_r_3__decode__me_nop_v_, calc_stage_r_3__decode__pipe_comp_v_, calc_stage_r_3__decode__pipe_int_v_, calc_stage_r_3__decode__pipe_mul_v_, calc_stage_r_3__decode__pipe_mem_v_, calc_stage_r_3__decode__pipe_fp_v_, calc_stage_r_3__decode__irf_w_v_, calc_stage_r_3__decode__frf_w_v_, calc_stage_r_3__decode__mhartid_r_v_, calc_stage_r_3__decode__dcache_w_v_, calc_stage_r_3__decode__dcache_r_v_, calc_stage_r_3__decode__fp_not_int_v_, calc_stage_r_3__decode__ret_v_, calc_stage_r_3__decode__amo_v_, calc_stage_r_3__decode__jmp_v_, calc_stage_r_3__decode__br_v_, calc_stage_r_3__decode__opw_v_, calc_stage_r_3__decode__fu_op__fu_op__3_, calc_stage_r_3__decode__fu_op__fu_op__2_, calc_stage_r_3__decode__fu_op__fu_op__1_, calc_stage_r_3__decode__fu_op__fu_op__0_, calc_stage_r_3__decode__rs1_addr__4_, calc_stage_r_3__decode__rs1_addr__3_, calc_stage_r_3__decode__rs1_addr__2_, calc_stage_r_3__decode__rs1_addr__1_, calc_stage_r_3__decode__rs1_addr__0_, calc_stage_r_3__decode__rs2_addr__4_, calc_stage_r_3__decode__rs2_addr__3_, calc_stage_r_3__decode__rs2_addr__2_, calc_stage_r_3__decode__rs2_addr__1_, calc_stage_r_3__decode__rs2_addr__0_, calc_status_o[103:99], calc_stage_r_3__decode__src1_sel_, calc_stage_r_3__decode__src2_sel_, calc_stage_r_3__decode__baddr_sel_, calc_stage_r_3__decode__result_sel_, calc_stage_r_2__instr_metadata__itag__7_, calc_stage_r_2__instr_metadata__itag__6_, calc_stage_r_2__instr_metadata__itag__5_, calc_stage_r_2__instr_metadata__itag__4_, calc_stage_r_2__instr_metadata__itag__3_, calc_stage_r_2__instr_metadata__itag__2_, calc_stage_r_2__instr_metadata__itag__1_, calc_stage_r_2__instr_metadata__itag__0_, calc_status_o[67:4], calc_stage_r_2__instr_metadata__fe_exception_not_instr_, calc_stage_r_2__instr_metadata__fe_exception_code__1_, calc_stage_r_2__instr_metadata__fe_exception_code__0_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__35_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__34_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__33_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__32_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__31_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__30_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__29_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__28_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__27_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__26_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__25_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__24_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__23_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__22_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__21_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__20_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__19_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__18_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__17_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__16_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__15_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__14_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__13_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__12_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__11_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__10_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__9_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__8_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__7_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__6_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__5_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__4_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__3_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__2_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__1_, calc_stage_r_2__instr_metadata__branch_metadata_fwd__0_, calc_stage_r_2__instr__31_, calc_stage_r_2__instr__30_, calc_stage_r_2__instr__29_, calc_stage_r_2__instr__28_, calc_stage_r_2__instr__27_, calc_stage_r_2__instr__26_, calc_stage_r_2__instr__25_, calc_stage_r_2__instr__24_, calc_stage_r_2__instr__23_, calc_stage_r_2__instr__22_, calc_stage_r_2__instr__21_, calc_stage_r_2__instr__20_, calc_stage_r_2__instr__19_, calc_stage_r_2__instr__18_, calc_stage_r_2__instr__17_, calc_stage_r_2__instr__16_, calc_stage_r_2__instr__15_, calc_stage_r_2__instr__14_, calc_stage_r_2__instr__13_, calc_stage_r_2__instr__12_, calc_stage_r_2__instr__11_, calc_stage_r_2__instr__10_, calc_stage_r_2__instr__9_, calc_stage_r_2__instr__8_, calc_stage_r_2__instr__7_, calc_stage_r_2__instr__6_, calc_stage_r_2__instr__5_, calc_stage_r_2__instr__4_, calc_stage_r_2__instr__3_, calc_stage_r_2__instr__2_, calc_stage_r_2__instr__1_, calc_stage_r_2__instr__0_, calc_stage_r_2__instr_operands__rs1__63_, calc_stage_r_2__instr_operands__rs1__62_, calc_stage_r_2__instr_operands__rs1__61_, calc_stage_r_2__instr_operands__rs1__60_, calc_stage_r_2__instr_operands__rs1__59_, calc_stage_r_2__instr_operands__rs1__58_, calc_stage_r_2__instr_operands__rs1__57_, calc_stage_r_2__instr_operands__rs1__56_, calc_stage_r_2__instr_operands__rs1__55_, calc_stage_r_2__instr_operands__rs1__54_, calc_stage_r_2__instr_operands__rs1__53_, calc_stage_r_2__instr_operands__rs1__52_, calc_stage_r_2__instr_operands__rs1__51_, calc_stage_r_2__instr_operands__rs1__50_, calc_stage_r_2__instr_operands__rs1__49_, calc_stage_r_2__instr_operands__rs1__48_, calc_stage_r_2__instr_operands__rs1__47_, calc_stage_r_2__instr_operands__rs1__46_, calc_stage_r_2__instr_operands__rs1__45_, calc_stage_r_2__instr_operands__rs1__44_, calc_stage_r_2__instr_operands__rs1__43_, calc_stage_r_2__instr_operands__rs1__42_, calc_stage_r_2__instr_operands__rs1__41_, calc_stage_r_2__instr_operands__rs1__40_, calc_stage_r_2__instr_operands__rs1__39_, calc_stage_r_2__instr_operands__rs1__38_, calc_stage_r_2__instr_operands__rs1__37_, calc_stage_r_2__instr_operands__rs1__36_, calc_stage_r_2__instr_operands__rs1__35_, calc_stage_r_2__instr_operands__rs1__34_, calc_stage_r_2__instr_operands__rs1__33_, calc_stage_r_2__instr_operands__rs1__32_, calc_stage_r_2__instr_operands__rs1__31_, calc_stage_r_2__instr_operands__rs1__30_, calc_stage_r_2__instr_operands__rs1__29_, calc_stage_r_2__instr_operands__rs1__28_, calc_stage_r_2__instr_operands__rs1__27_, calc_stage_r_2__instr_operands__rs1__26_, calc_stage_r_2__instr_operands__rs1__25_, calc_stage_r_2__instr_operands__rs1__24_, calc_stage_r_2__instr_operands__rs1__23_, calc_stage_r_2__instr_operands__rs1__22_, calc_stage_r_2__instr_operands__rs1__21_, calc_stage_r_2__instr_operands__rs1__20_, calc_stage_r_2__instr_operands__rs1__19_, calc_stage_r_2__instr_operands__rs1__18_, calc_stage_r_2__instr_operands__rs1__17_, calc_stage_r_2__instr_operands__rs1__16_, calc_stage_r_2__instr_operands__rs1__15_, calc_stage_r_2__instr_operands__rs1__14_, calc_stage_r_2__instr_operands__rs1__13_, calc_stage_r_2__instr_operands__rs1__12_, calc_stage_r_2__instr_operands__rs1__11_, calc_stage_r_2__instr_operands__rs1__10_, calc_stage_r_2__instr_operands__rs1__9_, calc_stage_r_2__instr_operands__rs1__8_, calc_stage_r_2__instr_operands__rs1__7_, calc_stage_r_2__instr_operands__rs1__6_, calc_stage_r_2__instr_operands__rs1__5_, calc_stage_r_2__instr_operands__rs1__4_, calc_stage_r_2__instr_operands__rs1__3_, calc_stage_r_2__instr_operands__rs1__2_, calc_stage_r_2__instr_operands__rs1__1_, calc_stage_r_2__instr_operands__rs1__0_, calc_stage_r_2__instr_operands__rs2__63_, calc_stage_r_2__instr_operands__rs2__62_, calc_stage_r_2__instr_operands__rs2__61_, calc_stage_r_2__instr_operands__rs2__60_, calc_stage_r_2__instr_operands__rs2__59_, calc_stage_r_2__instr_operands__rs2__58_, calc_stage_r_2__instr_operands__rs2__57_, calc_stage_r_2__instr_operands__rs2__56_, calc_stage_r_2__instr_operands__rs2__55_, calc_stage_r_2__instr_operands__rs2__54_, calc_stage_r_2__instr_operands__rs2__53_, calc_stage_r_2__instr_operands__rs2__52_, calc_stage_r_2__instr_operands__rs2__51_, calc_stage_r_2__instr_operands__rs2__50_, calc_stage_r_2__instr_operands__rs2__49_, calc_stage_r_2__instr_operands__rs2__48_, calc_stage_r_2__instr_operands__rs2__47_, calc_stage_r_2__instr_operands__rs2__46_, calc_stage_r_2__instr_operands__rs2__45_, calc_stage_r_2__instr_operands__rs2__44_, calc_stage_r_2__instr_operands__rs2__43_, calc_stage_r_2__instr_operands__rs2__42_, calc_stage_r_2__instr_operands__rs2__41_, calc_stage_r_2__instr_operands__rs2__40_, calc_stage_r_2__instr_operands__rs2__39_, calc_stage_r_2__instr_operands__rs2__38_, calc_stage_r_2__instr_operands__rs2__37_, calc_stage_r_2__instr_operands__rs2__36_, calc_stage_r_2__instr_operands__rs2__35_, calc_stage_r_2__instr_operands__rs2__34_, calc_stage_r_2__instr_operands__rs2__33_, calc_stage_r_2__instr_operands__rs2__32_, calc_stage_r_2__instr_operands__rs2__31_, calc_stage_r_2__instr_operands__rs2__30_, calc_stage_r_2__instr_operands__rs2__29_, calc_stage_r_2__instr_operands__rs2__28_, calc_stage_r_2__instr_operands__rs2__27_, calc_stage_r_2__instr_operands__rs2__26_, calc_stage_r_2__instr_operands__rs2__25_, calc_stage_r_2__instr_operands__rs2__24_, calc_stage_r_2__instr_operands__rs2__23_, calc_stage_r_2__instr_operands__rs2__22_, calc_stage_r_2__instr_operands__rs2__21_, calc_stage_r_2__instr_operands__rs2__20_, calc_stage_r_2__instr_operands__rs2__19_, calc_stage_r_2__instr_operands__rs2__18_, calc_stage_r_2__instr_operands__rs2__17_, calc_stage_r_2__instr_operands__rs2__16_, calc_stage_r_2__instr_operands__rs2__15_, calc_stage_r_2__instr_operands__rs2__14_, calc_stage_r_2__instr_operands__rs2__13_, calc_stage_r_2__instr_operands__rs2__12_, calc_stage_r_2__instr_operands__rs2__11_, calc_stage_r_2__instr_operands__rs2__10_, calc_stage_r_2__instr_operands__rs2__9_, calc_stage_r_2__instr_operands__rs2__8_, calc_stage_r_2__instr_operands__rs2__7_, calc_stage_r_2__instr_operands__rs2__6_, calc_stage_r_2__instr_operands__rs2__5_, calc_stage_r_2__instr_operands__rs2__4_, calc_stage_r_2__instr_operands__rs2__3_, calc_stage_r_2__instr_operands__rs2__2_, calc_stage_r_2__instr_operands__rs2__1_, calc_stage_r_2__instr_operands__rs2__0_, calc_stage_r_2__instr_operands__imm__63_, calc_stage_r_2__instr_operands__imm__62_, calc_stage_r_2__instr_operands__imm__61_, calc_stage_r_2__instr_operands__imm__60_, calc_stage_r_2__instr_operands__imm__59_, calc_stage_r_2__instr_operands__imm__58_, calc_stage_r_2__instr_operands__imm__57_, calc_stage_r_2__instr_operands__imm__56_, calc_stage_r_2__instr_operands__imm__55_, calc_stage_r_2__instr_operands__imm__54_, calc_stage_r_2__instr_operands__imm__53_, calc_stage_r_2__instr_operands__imm__52_, calc_stage_r_2__instr_operands__imm__51_, calc_stage_r_2__instr_operands__imm__50_, calc_stage_r_2__instr_operands__imm__49_, calc_stage_r_2__instr_operands__imm__48_, calc_stage_r_2__instr_operands__imm__47_, calc_stage_r_2__instr_operands__imm__46_, calc_stage_r_2__instr_operands__imm__45_, calc_stage_r_2__instr_operands__imm__44_, calc_stage_r_2__instr_operands__imm__43_, calc_stage_r_2__instr_operands__imm__42_, calc_stage_r_2__instr_operands__imm__41_, calc_stage_r_2__instr_operands__imm__40_, calc_stage_r_2__instr_operands__imm__39_, calc_stage_r_2__instr_operands__imm__38_, calc_stage_r_2__instr_operands__imm__37_, calc_stage_r_2__instr_operands__imm__36_, calc_stage_r_2__instr_operands__imm__35_, calc_stage_r_2__instr_operands__imm__34_, calc_stage_r_2__instr_operands__imm__33_, calc_stage_r_2__instr_operands__imm__32_, calc_stage_r_2__instr_operands__imm__31_, calc_stage_r_2__instr_operands__imm__30_, calc_stage_r_2__instr_operands__imm__29_, calc_stage_r_2__instr_operands__imm__28_, calc_stage_r_2__instr_operands__imm__27_, calc_stage_r_2__instr_operands__imm__26_, calc_stage_r_2__instr_operands__imm__25_, calc_stage_r_2__instr_operands__imm__24_, calc_stage_r_2__instr_operands__imm__23_, calc_stage_r_2__instr_operands__imm__22_, calc_stage_r_2__instr_operands__imm__21_, calc_stage_r_2__instr_operands__imm__20_, calc_stage_r_2__instr_operands__imm__19_, calc_stage_r_2__instr_operands__imm__18_, calc_stage_r_2__instr_operands__imm__17_, calc_stage_r_2__instr_operands__imm__16_, calc_stage_r_2__instr_operands__imm__15_, calc_stage_r_2__instr_operands__imm__14_, calc_stage_r_2__instr_operands__imm__13_, calc_stage_r_2__instr_operands__imm__12_, calc_stage_r_2__instr_operands__imm__11_, calc_stage_r_2__instr_operands__imm__10_, calc_stage_r_2__instr_operands__imm__9_, calc_stage_r_2__instr_operands__imm__8_, calc_stage_r_2__instr_operands__imm__7_, calc_stage_r_2__instr_operands__imm__6_, calc_stage_r_2__instr_operands__imm__5_, calc_stage_r_2__instr_operands__imm__4_, calc_stage_r_2__instr_operands__imm__3_, calc_stage_r_2__instr_operands__imm__2_, calc_stage_r_2__instr_operands__imm__1_, calc_stage_r_2__instr_operands__imm__0_, calc_stage_r_2__decode__instr_v_, calc_stage_r_2__decode__fe_nop_v_, calc_stage_r_2__decode__be_nop_v_, calc_stage_r_2__decode__me_nop_v_, calc_stage_r_2__decode__pipe_comp_v_, calc_stage_r_2__decode__pipe_int_v_, calc_stage_r_2__decode__pipe_mul_v_, calc_stage_r_2__decode__pipe_mem_v_, calc_stage_r_2__decode__pipe_fp_v_, calc_stage_r_2__decode__irf_w_v_, calc_stage_r_2__decode__frf_w_v_, calc_stage_r_2__decode__mhartid_r_v_, calc_stage_r_2__decode__dcache_w_v_, calc_stage_r_2__decode__dcache_r_v_, calc_stage_r_2__decode__fp_not_int_v_, calc_status_o[1:1], calc_stage_r_2__decode__amo_v_, calc_stage_r_2__decode__jmp_v_, calc_stage_r_2__decode__br_v_, calc_stage_r_2__decode__opw_v_, calc_stage_r_2__decode__fu_op__fu_op__3_, calc_stage_r_2__decode__fu_op__fu_op__2_, calc_stage_r_2__decode__fu_op__fu_op__1_, calc_stage_r_2__decode__fu_op__fu_op__0_, calc_stage_r_2__decode__rs1_addr__4_, calc_stage_r_2__decode__rs1_addr__3_, calc_stage_r_2__decode__rs1_addr__2_, calc_stage_r_2__decode__rs1_addr__1_, calc_stage_r_2__decode__rs1_addr__0_, calc_stage_r_2__decode__rs2_addr__4_, calc_stage_r_2__decode__rs2_addr__3_, calc_stage_r_2__decode__rs2_addr__2_, calc_stage_r_2__decode__rs2_addr__1_, calc_stage_r_2__decode__rs2_addr__0_, calc_status_o[93:89], calc_stage_r_2__decode__src1_sel_, calc_stage_r_2__decode__src2_sel_, calc_stage_r_2__decode__baddr_sel_, calc_stage_r_2__decode__result_sel_, calc_stage_r_1__instr_metadata__itag__7_, calc_stage_r_1__instr_metadata__itag__6_, calc_stage_r_1__instr_metadata__itag__5_, calc_stage_r_1__instr_metadata__itag__4_, calc_stage_r_1__instr_metadata__itag__3_, calc_stage_r_1__instr_metadata__itag__2_, calc_stage_r_1__instr_metadata__itag__1_, calc_stage_r_1__instr_metadata__itag__0_, calc_stage_r_1__instr_metadata__pc__63_, calc_stage_r_1__instr_metadata__pc__62_, calc_stage_r_1__instr_metadata__pc__61_, calc_stage_r_1__instr_metadata__pc__60_, calc_stage_r_1__instr_metadata__pc__59_, calc_stage_r_1__instr_metadata__pc__58_, calc_stage_r_1__instr_metadata__pc__57_, calc_stage_r_1__instr_metadata__pc__56_, calc_stage_r_1__instr_metadata__pc__55_, calc_stage_r_1__instr_metadata__pc__54_, calc_stage_r_1__instr_metadata__pc__53_, calc_stage_r_1__instr_metadata__pc__52_, calc_stage_r_1__instr_metadata__pc__51_, calc_stage_r_1__instr_metadata__pc__50_, calc_stage_r_1__instr_metadata__pc__49_, calc_stage_r_1__instr_metadata__pc__48_, calc_stage_r_1__instr_metadata__pc__47_, calc_stage_r_1__instr_metadata__pc__46_, calc_stage_r_1__instr_metadata__pc__45_, calc_stage_r_1__instr_metadata__pc__44_, calc_stage_r_1__instr_metadata__pc__43_, calc_stage_r_1__instr_metadata__pc__42_, calc_stage_r_1__instr_metadata__pc__41_, calc_stage_r_1__instr_metadata__pc__40_, calc_stage_r_1__instr_metadata__pc__39_, calc_stage_r_1__instr_metadata__pc__38_, calc_stage_r_1__instr_metadata__pc__37_, calc_stage_r_1__instr_metadata__pc__36_, calc_stage_r_1__instr_metadata__pc__35_, calc_stage_r_1__instr_metadata__pc__34_, calc_stage_r_1__instr_metadata__pc__33_, calc_stage_r_1__instr_metadata__pc__32_, calc_stage_r_1__instr_metadata__pc__31_, calc_stage_r_1__instr_metadata__pc__30_, calc_stage_r_1__instr_metadata__pc__29_, calc_stage_r_1__instr_metadata__pc__28_, calc_stage_r_1__instr_metadata__pc__27_, calc_stage_r_1__instr_metadata__pc__26_, calc_stage_r_1__instr_metadata__pc__25_, calc_stage_r_1__instr_metadata__pc__24_, calc_stage_r_1__instr_metadata__pc__23_, calc_stage_r_1__instr_metadata__pc__22_, calc_stage_r_1__instr_metadata__pc__21_, calc_stage_r_1__instr_metadata__pc__20_, calc_stage_r_1__instr_metadata__pc__19_, calc_stage_r_1__instr_metadata__pc__18_, calc_stage_r_1__instr_metadata__pc__17_, calc_stage_r_1__instr_metadata__pc__16_, calc_stage_r_1__instr_metadata__pc__15_, calc_stage_r_1__instr_metadata__pc__14_, calc_stage_r_1__instr_metadata__pc__13_, calc_stage_r_1__instr_metadata__pc__12_, calc_stage_r_1__instr_metadata__pc__11_, calc_stage_r_1__instr_metadata__pc__10_, calc_stage_r_1__instr_metadata__pc__9_, calc_stage_r_1__instr_metadata__pc__8_, calc_stage_r_1__instr_metadata__pc__7_, calc_stage_r_1__instr_metadata__pc__6_, calc_stage_r_1__instr_metadata__pc__5_, calc_stage_r_1__instr_metadata__pc__4_, calc_stage_r_1__instr_metadata__pc__3_, calc_stage_r_1__instr_metadata__pc__2_, calc_stage_r_1__instr_metadata__pc__1_, calc_stage_r_1__instr_metadata__pc__0_, calc_stage_r_1__instr_metadata__fe_exception_not_instr_, calc_stage_r_1__instr_metadata__fe_exception_code__1_, calc_stage_r_1__instr_metadata__fe_exception_code__0_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__35_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__34_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__33_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__32_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__31_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__30_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__29_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__28_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__27_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__26_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__25_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__24_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__23_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__22_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__21_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__20_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__19_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__18_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__17_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__16_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__15_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__14_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__13_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__12_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__11_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__10_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__9_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__8_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__7_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__6_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__5_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__4_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__3_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__2_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__1_, calc_stage_r_1__instr_metadata__branch_metadata_fwd__0_, calc_stage_r_1__instr__31_, calc_stage_r_1__instr__30_, calc_stage_r_1__instr__29_, calc_stage_r_1__instr__28_, calc_stage_r_1__instr__27_, calc_stage_r_1__instr__26_, calc_stage_r_1__instr__25_, calc_stage_r_1__instr__24_, calc_stage_r_1__instr__23_, calc_stage_r_1__instr__22_, calc_stage_r_1__instr__21_, calc_stage_r_1__instr__20_, calc_stage_r_1__instr__19_, calc_stage_r_1__instr__18_, calc_stage_r_1__instr__17_, calc_stage_r_1__instr__16_, calc_stage_r_1__instr__15_, calc_stage_r_1__instr__14_, calc_stage_r_1__instr__13_, calc_stage_r_1__instr__12_, calc_stage_r_1__instr__11_, calc_stage_r_1__instr__10_, calc_stage_r_1__instr__9_, calc_stage_r_1__instr__8_, calc_stage_r_1__instr__7_, calc_stage_r_1__instr__6_, calc_stage_r_1__instr__5_, calc_stage_r_1__instr__4_, calc_stage_r_1__instr__3_, calc_stage_r_1__instr__2_, calc_stage_r_1__instr__1_, calc_stage_r_1__instr__0_, calc_stage_r_1__instr_operands__rs1__63_, calc_stage_r_1__instr_operands__rs1__62_, calc_stage_r_1__instr_operands__rs1__61_, calc_stage_r_1__instr_operands__rs1__60_, calc_stage_r_1__instr_operands__rs1__59_, calc_stage_r_1__instr_operands__rs1__58_, calc_stage_r_1__instr_operands__rs1__57_, calc_stage_r_1__instr_operands__rs1__56_, calc_stage_r_1__instr_operands__rs1__55_, calc_stage_r_1__instr_operands__rs1__54_, calc_stage_r_1__instr_operands__rs1__53_, calc_stage_r_1__instr_operands__rs1__52_, calc_stage_r_1__instr_operands__rs1__51_, calc_stage_r_1__instr_operands__rs1__50_, calc_stage_r_1__instr_operands__rs1__49_, calc_stage_r_1__instr_operands__rs1__48_, calc_stage_r_1__instr_operands__rs1__47_, calc_stage_r_1__instr_operands__rs1__46_, calc_stage_r_1__instr_operands__rs1__45_, calc_stage_r_1__instr_operands__rs1__44_, calc_stage_r_1__instr_operands__rs1__43_, calc_stage_r_1__instr_operands__rs1__42_, calc_stage_r_1__instr_operands__rs1__41_, calc_stage_r_1__instr_operands__rs1__40_, calc_stage_r_1__instr_operands__rs1__39_, calc_stage_r_1__instr_operands__rs1__38_, calc_stage_r_1__instr_operands__rs1__37_, calc_stage_r_1__instr_operands__rs1__36_, calc_stage_r_1__instr_operands__rs1__35_, calc_stage_r_1__instr_operands__rs1__34_, calc_stage_r_1__instr_operands__rs1__33_, calc_stage_r_1__instr_operands__rs1__32_, calc_stage_r_1__instr_operands__rs1__31_, calc_stage_r_1__instr_operands__rs1__30_, calc_stage_r_1__instr_operands__rs1__29_, calc_stage_r_1__instr_operands__rs1__28_, calc_stage_r_1__instr_operands__rs1__27_, calc_stage_r_1__instr_operands__rs1__26_, calc_stage_r_1__instr_operands__rs1__25_, calc_stage_r_1__instr_operands__rs1__24_, calc_stage_r_1__instr_operands__rs1__23_, calc_stage_r_1__instr_operands__rs1__22_, calc_stage_r_1__instr_operands__rs1__21_, calc_stage_r_1__instr_operands__rs1__20_, calc_stage_r_1__instr_operands__rs1__19_, calc_stage_r_1__instr_operands__rs1__18_, calc_stage_r_1__instr_operands__rs1__17_, calc_stage_r_1__instr_operands__rs1__16_, calc_stage_r_1__instr_operands__rs1__15_, calc_stage_r_1__instr_operands__rs1__14_, calc_stage_r_1__instr_operands__rs1__13_, calc_stage_r_1__instr_operands__rs1__12_, calc_stage_r_1__instr_operands__rs1__11_, calc_stage_r_1__instr_operands__rs1__10_, calc_stage_r_1__instr_operands__rs1__9_, calc_stage_r_1__instr_operands__rs1__8_, calc_stage_r_1__instr_operands__rs1__7_, calc_stage_r_1__instr_operands__rs1__6_, calc_stage_r_1__instr_operands__rs1__5_, calc_stage_r_1__instr_operands__rs1__4_, calc_stage_r_1__instr_operands__rs1__3_, calc_stage_r_1__instr_operands__rs1__2_, calc_stage_r_1__instr_operands__rs1__1_, calc_stage_r_1__instr_operands__rs1__0_, calc_stage_r_1__instr_operands__rs2__63_, calc_stage_r_1__instr_operands__rs2__62_, calc_stage_r_1__instr_operands__rs2__61_, calc_stage_r_1__instr_operands__rs2__60_, calc_stage_r_1__instr_operands__rs2__59_, calc_stage_r_1__instr_operands__rs2__58_, calc_stage_r_1__instr_operands__rs2__57_, calc_stage_r_1__instr_operands__rs2__56_, calc_stage_r_1__instr_operands__rs2__55_, calc_stage_r_1__instr_operands__rs2__54_, calc_stage_r_1__instr_operands__rs2__53_, calc_stage_r_1__instr_operands__rs2__52_, calc_stage_r_1__instr_operands__rs2__51_, calc_stage_r_1__instr_operands__rs2__50_, calc_stage_r_1__instr_operands__rs2__49_, calc_stage_r_1__instr_operands__rs2__48_, calc_stage_r_1__instr_operands__rs2__47_, calc_stage_r_1__instr_operands__rs2__46_, calc_stage_r_1__instr_operands__rs2__45_, calc_stage_r_1__instr_operands__rs2__44_, calc_stage_r_1__instr_operands__rs2__43_, calc_stage_r_1__instr_operands__rs2__42_, calc_stage_r_1__instr_operands__rs2__41_, calc_stage_r_1__instr_operands__rs2__40_, calc_stage_r_1__instr_operands__rs2__39_, calc_stage_r_1__instr_operands__rs2__38_, calc_stage_r_1__instr_operands__rs2__37_, calc_stage_r_1__instr_operands__rs2__36_, calc_stage_r_1__instr_operands__rs2__35_, calc_stage_r_1__instr_operands__rs2__34_, calc_stage_r_1__instr_operands__rs2__33_, calc_stage_r_1__instr_operands__rs2__32_, calc_stage_r_1__instr_operands__rs2__31_, calc_stage_r_1__instr_operands__rs2__30_, calc_stage_r_1__instr_operands__rs2__29_, calc_stage_r_1__instr_operands__rs2__28_, calc_stage_r_1__instr_operands__rs2__27_, calc_stage_r_1__instr_operands__rs2__26_, calc_stage_r_1__instr_operands__rs2__25_, calc_stage_r_1__instr_operands__rs2__24_, calc_stage_r_1__instr_operands__rs2__23_, calc_stage_r_1__instr_operands__rs2__22_, calc_stage_r_1__instr_operands__rs2__21_, calc_stage_r_1__instr_operands__rs2__20_, calc_stage_r_1__instr_operands__rs2__19_, calc_stage_r_1__instr_operands__rs2__18_, calc_stage_r_1__instr_operands__rs2__17_, calc_stage_r_1__instr_operands__rs2__16_, calc_stage_r_1__instr_operands__rs2__15_, calc_stage_r_1__instr_operands__rs2__14_, calc_stage_r_1__instr_operands__rs2__13_, calc_stage_r_1__instr_operands__rs2__12_, calc_stage_r_1__instr_operands__rs2__11_, calc_stage_r_1__instr_operands__rs2__10_, calc_stage_r_1__instr_operands__rs2__9_, calc_stage_r_1__instr_operands__rs2__8_, calc_stage_r_1__instr_operands__rs2__7_, calc_stage_r_1__instr_operands__rs2__6_, calc_stage_r_1__instr_operands__rs2__5_, calc_stage_r_1__instr_operands__rs2__4_, calc_stage_r_1__instr_operands__rs2__3_, calc_stage_r_1__instr_operands__rs2__2_, calc_stage_r_1__instr_operands__rs2__1_, calc_stage_r_1__instr_operands__rs2__0_, calc_stage_r_1__instr_operands__imm__63_, calc_stage_r_1__instr_operands__imm__62_, calc_stage_r_1__instr_operands__imm__61_, calc_stage_r_1__instr_operands__imm__60_, calc_stage_r_1__instr_operands__imm__59_, calc_stage_r_1__instr_operands__imm__58_, calc_stage_r_1__instr_operands__imm__57_, calc_stage_r_1__instr_operands__imm__56_, calc_stage_r_1__instr_operands__imm__55_, calc_stage_r_1__instr_operands__imm__54_, calc_stage_r_1__instr_operands__imm__53_, calc_stage_r_1__instr_operands__imm__52_, calc_stage_r_1__instr_operands__imm__51_, calc_stage_r_1__instr_operands__imm__50_, calc_stage_r_1__instr_operands__imm__49_, calc_stage_r_1__instr_operands__imm__48_, calc_stage_r_1__instr_operands__imm__47_, calc_stage_r_1__instr_operands__imm__46_, calc_stage_r_1__instr_operands__imm__45_, calc_stage_r_1__instr_operands__imm__44_, calc_stage_r_1__instr_operands__imm__43_, calc_stage_r_1__instr_operands__imm__42_, calc_stage_r_1__instr_operands__imm__41_, calc_stage_r_1__instr_operands__imm__40_, calc_stage_r_1__instr_operands__imm__39_, calc_stage_r_1__instr_operands__imm__38_, calc_stage_r_1__instr_operands__imm__37_, calc_stage_r_1__instr_operands__imm__36_, calc_stage_r_1__instr_operands__imm__35_, calc_stage_r_1__instr_operands__imm__34_, calc_stage_r_1__instr_operands__imm__33_, calc_stage_r_1__instr_operands__imm__32_, calc_stage_r_1__instr_operands__imm__31_, calc_stage_r_1__instr_operands__imm__30_, calc_stage_r_1__instr_operands__imm__29_, calc_stage_r_1__instr_operands__imm__28_, calc_stage_r_1__instr_operands__imm__27_, calc_stage_r_1__instr_operands__imm__26_, calc_stage_r_1__instr_operands__imm__25_, calc_stage_r_1__instr_operands__imm__24_, calc_stage_r_1__instr_operands__imm__23_, calc_stage_r_1__instr_operands__imm__22_, calc_stage_r_1__instr_operands__imm__21_, calc_stage_r_1__instr_operands__imm__20_, calc_stage_r_1__instr_operands__imm__19_, calc_stage_r_1__instr_operands__imm__18_, calc_stage_r_1__instr_operands__imm__17_, calc_stage_r_1__instr_operands__imm__16_, calc_stage_r_1__instr_operands__imm__15_, calc_stage_r_1__instr_operands__imm__14_, calc_stage_r_1__instr_operands__imm__13_, calc_stage_r_1__instr_operands__imm__12_, calc_stage_r_1__instr_operands__imm__11_, calc_stage_r_1__instr_operands__imm__10_, calc_stage_r_1__instr_operands__imm__9_, calc_stage_r_1__instr_operands__imm__8_, calc_stage_r_1__instr_operands__imm__7_, calc_stage_r_1__instr_operands__imm__6_, calc_stage_r_1__instr_operands__imm__5_, calc_stage_r_1__instr_operands__imm__4_, calc_stage_r_1__instr_operands__imm__3_, calc_stage_r_1__instr_operands__imm__2_, calc_stage_r_1__instr_operands__imm__1_, calc_stage_r_1__instr_operands__imm__0_, calc_stage_r_1__decode__instr_v_, calc_stage_r_1__decode__fe_nop_v_, calc_stage_r_1__decode__be_nop_v_, calc_stage_r_1__decode__me_nop_v_, calc_stage_r_1__decode__pipe_comp_v_, calc_stage_r_1__decode__pipe_int_v_, calc_stage_r_1__decode__pipe_mul_v_, calc_stage_r_1__decode__pipe_mem_v_, calc_stage_r_1__decode__pipe_fp_v_, calc_stage_r_1__decode__irf_w_v_, calc_stage_r_1__decode__frf_w_v_, calc_stage_r_1__decode__mhartid_r_v_, calc_stage_r_1__decode__dcache_w_v_, calc_stage_r_1__decode__dcache_r_v_, calc_stage_r_1__decode__fp_not_int_v_, calc_stage_r_1__decode__ret_v_, calc_stage_r_1__decode__amo_v_, calc_stage_r_1__decode__jmp_v_, calc_stage_r_1__decode__br_v_, calc_stage_r_1__decode__opw_v_, calc_stage_r_1__decode__fu_op__fu_op__3_, calc_stage_r_1__decode__fu_op__fu_op__2_, calc_stage_r_1__decode__fu_op__fu_op__1_, calc_stage_r_1__decode__fu_op__fu_op__0_, calc_stage_r_1__decode__rs1_addr__4_, calc_stage_r_1__decode__rs1_addr__3_, calc_stage_r_1__decode__rs1_addr__2_, calc_stage_r_1__decode__rs1_addr__1_, calc_stage_r_1__decode__rs1_addr__0_, calc_stage_r_1__decode__rs2_addr__4_, calc_stage_r_1__decode__rs2_addr__3_, calc_stage_r_1__decode__rs2_addr__2_, calc_stage_r_1__decode__rs2_addr__1_, calc_stage_r_1__decode__rs2_addr__0_, calc_status_o[83:79], calc_stage_r_1__decode__src1_sel_, calc_stage_r_1__decode__src2_sel_, calc_stage_r_1__decode__baddr_sel_, calc_stage_r_1__decode__result_sel_, calc_stage_r_0__instr_metadata__itag__7_, calc_stage_r_0__instr_metadata__itag__6_, calc_stage_r_0__instr_metadata__itag__5_, calc_stage_r_0__instr_metadata__itag__4_, calc_stage_r_0__instr_metadata__itag__3_, calc_stage_r_0__instr_metadata__itag__2_, calc_stage_r_0__instr_metadata__itag__1_, calc_stage_r_0__instr_metadata__itag__0_, calc_stage_r_0__instr_metadata__pc__63_, calc_stage_r_0__instr_metadata__pc__62_, calc_stage_r_0__instr_metadata__pc__61_, calc_stage_r_0__instr_metadata__pc__60_, calc_stage_r_0__instr_metadata__pc__59_, calc_stage_r_0__instr_metadata__pc__58_, calc_stage_r_0__instr_metadata__pc__57_, calc_stage_r_0__instr_metadata__pc__56_, calc_stage_r_0__instr_metadata__pc__55_, calc_stage_r_0__instr_metadata__pc__54_, calc_stage_r_0__instr_metadata__pc__53_, calc_stage_r_0__instr_metadata__pc__52_, calc_stage_r_0__instr_metadata__pc__51_, calc_stage_r_0__instr_metadata__pc__50_, calc_stage_r_0__instr_metadata__pc__49_, calc_stage_r_0__instr_metadata__pc__48_, calc_stage_r_0__instr_metadata__pc__47_, calc_stage_r_0__instr_metadata__pc__46_, calc_stage_r_0__instr_metadata__pc__45_, calc_stage_r_0__instr_metadata__pc__44_, calc_stage_r_0__instr_metadata__pc__43_, calc_stage_r_0__instr_metadata__pc__42_, calc_stage_r_0__instr_metadata__pc__41_, calc_stage_r_0__instr_metadata__pc__40_, calc_stage_r_0__instr_metadata__pc__39_, calc_stage_r_0__instr_metadata__pc__38_, calc_stage_r_0__instr_metadata__pc__37_, calc_stage_r_0__instr_metadata__pc__36_, calc_stage_r_0__instr_metadata__pc__35_, calc_stage_r_0__instr_metadata__pc__34_, calc_stage_r_0__instr_metadata__pc__33_, calc_stage_r_0__instr_metadata__pc__32_, calc_stage_r_0__instr_metadata__pc__31_, calc_stage_r_0__instr_metadata__pc__30_, calc_stage_r_0__instr_metadata__pc__29_, calc_stage_r_0__instr_metadata__pc__28_, calc_stage_r_0__instr_metadata__pc__27_, calc_stage_r_0__instr_metadata__pc__26_, calc_stage_r_0__instr_metadata__pc__25_, calc_stage_r_0__instr_metadata__pc__24_, calc_stage_r_0__instr_metadata__pc__23_, calc_stage_r_0__instr_metadata__pc__22_, calc_stage_r_0__instr_metadata__pc__21_, calc_stage_r_0__instr_metadata__pc__20_, calc_stage_r_0__instr_metadata__pc__19_, calc_stage_r_0__instr_metadata__pc__18_, calc_stage_r_0__instr_metadata__pc__17_, calc_stage_r_0__instr_metadata__pc__16_, calc_stage_r_0__instr_metadata__pc__15_, calc_stage_r_0__instr_metadata__pc__14_, calc_stage_r_0__instr_metadata__pc__13_, calc_stage_r_0__instr_metadata__pc__12_, calc_stage_r_0__instr_metadata__pc__11_, calc_stage_r_0__instr_metadata__pc__10_, calc_stage_r_0__instr_metadata__pc__9_, calc_stage_r_0__instr_metadata__pc__8_, calc_stage_r_0__instr_metadata__pc__7_, calc_stage_r_0__instr_metadata__pc__6_, calc_stage_r_0__instr_metadata__pc__5_, calc_stage_r_0__instr_metadata__pc__4_, calc_stage_r_0__instr_metadata__pc__3_, calc_stage_r_0__instr_metadata__pc__2_, calc_stage_r_0__instr_metadata__pc__1_, calc_stage_r_0__instr_metadata__pc__0_, calc_stage_r_0__instr_metadata__fe_exception_not_instr_, calc_stage_r_0__instr_metadata__fe_exception_code__1_, calc_stage_r_0__instr_metadata__fe_exception_code__0_, calc_status_o[157:122], calc_stage_r_0__instr__31_, calc_stage_r_0__instr__30_, calc_stage_r_0__instr__29_, calc_stage_r_0__instr__28_, calc_stage_r_0__instr__27_, calc_stage_r_0__instr__26_, calc_stage_r_0__instr__25_, calc_stage_r_0__instr__24_, calc_stage_r_0__instr__23_, calc_stage_r_0__instr__22_, calc_stage_r_0__instr__21_, calc_stage_r_0__instr__20_, calc_stage_r_0__instr__19_, calc_stage_r_0__instr__18_, calc_stage_r_0__instr__17_, calc_stage_r_0__instr__16_, calc_stage_r_0__instr__15_, calc_stage_r_0__instr__14_, calc_stage_r_0__instr__13_, calc_stage_r_0__instr__12_, calc_stage_r_0__instr__11_, calc_stage_r_0__instr__10_, calc_stage_r_0__instr__9_, calc_stage_r_0__instr__8_, calc_stage_r_0__instr__7_, calc_stage_r_0__instr__6_, calc_stage_r_0__instr__5_, calc_stage_r_0__instr__4_, calc_stage_r_0__instr__3_, calc_stage_r_0__instr__2_, calc_stage_r_0__instr__1_, calc_stage_r_0__instr__0_, calc_stage_r_0__instr_operands__rs1__63_, calc_stage_r_0__instr_operands__rs1__62_, calc_stage_r_0__instr_operands__rs1__61_, calc_stage_r_0__instr_operands__rs1__60_, calc_stage_r_0__instr_operands__rs1__59_, calc_stage_r_0__instr_operands__rs1__58_, calc_stage_r_0__instr_operands__rs1__57_, calc_stage_r_0__instr_operands__rs1__56_, calc_stage_r_0__instr_operands__rs1__55_, calc_stage_r_0__instr_operands__rs1__54_, calc_stage_r_0__instr_operands__rs1__53_, calc_stage_r_0__instr_operands__rs1__52_, calc_stage_r_0__instr_operands__rs1__51_, calc_stage_r_0__instr_operands__rs1__50_, calc_stage_r_0__instr_operands__rs1__49_, calc_stage_r_0__instr_operands__rs1__48_, calc_stage_r_0__instr_operands__rs1__47_, calc_stage_r_0__instr_operands__rs1__46_, calc_stage_r_0__instr_operands__rs1__45_, calc_stage_r_0__instr_operands__rs1__44_, calc_stage_r_0__instr_operands__rs1__43_, calc_stage_r_0__instr_operands__rs1__42_, calc_stage_r_0__instr_operands__rs1__41_, calc_stage_r_0__instr_operands__rs1__40_, calc_stage_r_0__instr_operands__rs1__39_, calc_stage_r_0__instr_operands__rs1__38_, calc_stage_r_0__instr_operands__rs1__37_, calc_stage_r_0__instr_operands__rs1__36_, calc_stage_r_0__instr_operands__rs1__35_, calc_stage_r_0__instr_operands__rs1__34_, calc_stage_r_0__instr_operands__rs1__33_, calc_stage_r_0__instr_operands__rs1__32_, calc_stage_r_0__instr_operands__rs1__31_, calc_stage_r_0__instr_operands__rs1__30_, calc_stage_r_0__instr_operands__rs1__29_, calc_stage_r_0__instr_operands__rs1__28_, calc_stage_r_0__instr_operands__rs1__27_, calc_stage_r_0__instr_operands__rs1__26_, calc_stage_r_0__instr_operands__rs1__25_, calc_stage_r_0__instr_operands__rs1__24_, calc_stage_r_0__instr_operands__rs1__23_, calc_stage_r_0__instr_operands__rs1__22_, calc_stage_r_0__instr_operands__rs1__21_, calc_stage_r_0__instr_operands__rs1__20_, calc_stage_r_0__instr_operands__rs1__19_, calc_stage_r_0__instr_operands__rs1__18_, calc_stage_r_0__instr_operands__rs1__17_, calc_stage_r_0__instr_operands__rs1__16_, calc_stage_r_0__instr_operands__rs1__15_, calc_stage_r_0__instr_operands__rs1__14_, calc_stage_r_0__instr_operands__rs1__13_, calc_stage_r_0__instr_operands__rs1__12_, calc_stage_r_0__instr_operands__rs1__11_, calc_stage_r_0__instr_operands__rs1__10_, calc_stage_r_0__instr_operands__rs1__9_, calc_stage_r_0__instr_operands__rs1__8_, calc_stage_r_0__instr_operands__rs1__7_, calc_stage_r_0__instr_operands__rs1__6_, calc_stage_r_0__instr_operands__rs1__5_, calc_stage_r_0__instr_operands__rs1__4_, calc_stage_r_0__instr_operands__rs1__3_, calc_stage_r_0__instr_operands__rs1__2_, calc_stage_r_0__instr_operands__rs1__1_, calc_stage_r_0__instr_operands__rs1__0_, calc_stage_r_0__instr_operands__rs2__63_, calc_stage_r_0__instr_operands__rs2__62_, calc_stage_r_0__instr_operands__rs2__61_, calc_stage_r_0__instr_operands__rs2__60_, calc_stage_r_0__instr_operands__rs2__59_, calc_stage_r_0__instr_operands__rs2__58_, calc_stage_r_0__instr_operands__rs2__57_, calc_stage_r_0__instr_operands__rs2__56_, calc_stage_r_0__instr_operands__rs2__55_, calc_stage_r_0__instr_operands__rs2__54_, calc_stage_r_0__instr_operands__rs2__53_, calc_stage_r_0__instr_operands__rs2__52_, calc_stage_r_0__instr_operands__rs2__51_, calc_stage_r_0__instr_operands__rs2__50_, calc_stage_r_0__instr_operands__rs2__49_, calc_stage_r_0__instr_operands__rs2__48_, calc_stage_r_0__instr_operands__rs2__47_, calc_stage_r_0__instr_operands__rs2__46_, calc_stage_r_0__instr_operands__rs2__45_, calc_stage_r_0__instr_operands__rs2__44_, calc_stage_r_0__instr_operands__rs2__43_, calc_stage_r_0__instr_operands__rs2__42_, calc_stage_r_0__instr_operands__rs2__41_, calc_stage_r_0__instr_operands__rs2__40_, calc_stage_r_0__instr_operands__rs2__39_, calc_stage_r_0__instr_operands__rs2__38_, calc_stage_r_0__instr_operands__rs2__37_, calc_stage_r_0__instr_operands__rs2__36_, calc_stage_r_0__instr_operands__rs2__35_, calc_stage_r_0__instr_operands__rs2__34_, calc_stage_r_0__instr_operands__rs2__33_, calc_stage_r_0__instr_operands__rs2__32_, calc_stage_r_0__instr_operands__rs2__31_, calc_stage_r_0__instr_operands__rs2__30_, calc_stage_r_0__instr_operands__rs2__29_, calc_stage_r_0__instr_operands__rs2__28_, calc_stage_r_0__instr_operands__rs2__27_, calc_stage_r_0__instr_operands__rs2__26_, calc_stage_r_0__instr_operands__rs2__25_, calc_stage_r_0__instr_operands__rs2__24_, calc_stage_r_0__instr_operands__rs2__23_, calc_stage_r_0__instr_operands__rs2__22_, calc_stage_r_0__instr_operands__rs2__21_, calc_stage_r_0__instr_operands__rs2__20_, calc_stage_r_0__instr_operands__rs2__19_, calc_stage_r_0__instr_operands__rs2__18_, calc_stage_r_0__instr_operands__rs2__17_, calc_stage_r_0__instr_operands__rs2__16_, calc_stage_r_0__instr_operands__rs2__15_, calc_stage_r_0__instr_operands__rs2__14_, calc_stage_r_0__instr_operands__rs2__13_, calc_stage_r_0__instr_operands__rs2__12_, calc_stage_r_0__instr_operands__rs2__11_, calc_stage_r_0__instr_operands__rs2__10_, calc_stage_r_0__instr_operands__rs2__9_, calc_stage_r_0__instr_operands__rs2__8_, calc_stage_r_0__instr_operands__rs2__7_, calc_stage_r_0__instr_operands__rs2__6_, calc_stage_r_0__instr_operands__rs2__5_, calc_stage_r_0__instr_operands__rs2__4_, calc_stage_r_0__instr_operands__rs2__3_, calc_stage_r_0__instr_operands__rs2__2_, calc_stage_r_0__instr_operands__rs2__1_, calc_stage_r_0__instr_operands__rs2__0_, calc_stage_r_0__instr_operands__imm__63_, calc_stage_r_0__instr_operands__imm__62_, calc_stage_r_0__instr_operands__imm__61_, calc_stage_r_0__instr_operands__imm__60_, calc_stage_r_0__instr_operands__imm__59_, calc_stage_r_0__instr_operands__imm__58_, calc_stage_r_0__instr_operands__imm__57_, calc_stage_r_0__instr_operands__imm__56_, calc_stage_r_0__instr_operands__imm__55_, calc_stage_r_0__instr_operands__imm__54_, calc_stage_r_0__instr_operands__imm__53_, calc_stage_r_0__instr_operands__imm__52_, calc_stage_r_0__instr_operands__imm__51_, calc_stage_r_0__instr_operands__imm__50_, calc_stage_r_0__instr_operands__imm__49_, calc_stage_r_0__instr_operands__imm__48_, calc_stage_r_0__instr_operands__imm__47_, calc_stage_r_0__instr_operands__imm__46_, calc_stage_r_0__instr_operands__imm__45_, calc_stage_r_0__instr_operands__imm__44_, calc_stage_r_0__instr_operands__imm__43_, calc_stage_r_0__instr_operands__imm__42_, calc_stage_r_0__instr_operands__imm__41_, calc_stage_r_0__instr_operands__imm__40_, calc_stage_r_0__instr_operands__imm__39_, calc_stage_r_0__instr_operands__imm__38_, calc_stage_r_0__instr_operands__imm__37_, calc_stage_r_0__instr_operands__imm__36_, calc_stage_r_0__instr_operands__imm__35_, calc_stage_r_0__instr_operands__imm__34_, calc_stage_r_0__instr_operands__imm__33_, calc_stage_r_0__instr_operands__imm__32_, calc_stage_r_0__instr_operands__imm__31_, calc_stage_r_0__instr_operands__imm__30_, calc_stage_r_0__instr_operands__imm__29_, calc_stage_r_0__instr_operands__imm__28_, calc_stage_r_0__instr_operands__imm__27_, calc_stage_r_0__instr_operands__imm__26_, calc_stage_r_0__instr_operands__imm__25_, calc_stage_r_0__instr_operands__imm__24_, calc_stage_r_0__instr_operands__imm__23_, calc_stage_r_0__instr_operands__imm__22_, calc_stage_r_0__instr_operands__imm__21_, calc_stage_r_0__instr_operands__imm__20_, calc_stage_r_0__instr_operands__imm__19_, calc_stage_r_0__instr_operands__imm__18_, calc_stage_r_0__instr_operands__imm__17_, calc_stage_r_0__instr_operands__imm__16_, calc_stage_r_0__instr_operands__imm__15_, calc_stage_r_0__instr_operands__imm__14_, calc_stage_r_0__instr_operands__imm__13_, calc_stage_r_0__instr_operands__imm__12_, calc_stage_r_0__instr_operands__imm__11_, calc_stage_r_0__instr_operands__imm__10_, calc_stage_r_0__instr_operands__imm__9_, calc_stage_r_0__instr_operands__imm__8_, calc_stage_r_0__instr_operands__imm__7_, calc_stage_r_0__instr_operands__imm__6_, calc_stage_r_0__instr_operands__imm__5_, calc_stage_r_0__instr_operands__imm__4_, calc_stage_r_0__instr_operands__imm__3_, calc_stage_r_0__instr_operands__imm__2_, calc_stage_r_0__instr_operands__imm__1_, calc_stage_r_0__instr_operands__imm__0_, calc_stage_r_0__decode__instr_v_, calc_stage_r_0__decode__fe_nop_v_, calc_stage_r_0__decode__be_nop_v_, calc_stage_r_0__decode__me_nop_v_, calc_stage_r_0__decode__pipe_comp_v_, calc_stage_r_0__decode__pipe_int_v_, calc_stage_r_0__decode__pipe_mul_v_, calc_stage_r_0__decode__pipe_mem_v_, calc_stage_r_0__decode__pipe_fp_v_, calc_stage_r_0__decode__irf_w_v_, calc_stage_r_0__decode__frf_w_v_, calc_stage_r_0__decode__mhartid_r_v_, calc_stage_r_0__decode__dcache_w_v_, calc_stage_r_0__decode__dcache_r_v_, calc_stage_r_0__decode__fp_not_int_v_, calc_stage_r_0__decode__ret_v_, calc_stage_r_0__decode__amo_v_, calc_stage_r_0__decode__jmp_v_, calc_stage_r_0__decode__br_v_, calc_stage_r_0__decode__opw_v_, calc_stage_r_0__decode__fu_op__fu_op__3_, calc_stage_r_0__decode__fu_op__fu_op__2_, calc_stage_r_0__decode__fu_op__fu_op__1_, calc_stage_r_0__decode__fu_op__fu_op__0_, calc_stage_r_0__decode__rs1_addr__4_, calc_stage_r_0__decode__rs1_addr__3_, calc_stage_r_0__decode__rs1_addr__2_, calc_stage_r_0__decode__rs1_addr__1_, calc_stage_r_0__decode__rs1_addr__0_, calc_stage_r_0__decode__rs2_addr__4_, calc_stage_r_0__decode__rs2_addr__3_, calc_stage_r_0__decode__rs2_addr__2_, calc_stage_r_0__decode__rs2_addr__1_, calc_stage_r_0__decode__rs2_addr__0_, calc_status_o[73:69], calc_stage_r_0__decode__src1_sel_, calc_stage_r_0__decode__src2_sel_, calc_stage_r_0__decode__baddr_sel_, calc_stage_r_0__decode__result_sel_ })
  );


  bsg_mux_segmented_segments_p5_segment_width_p128
  comp_stage_mux
  (
    .data0_i({ comp_stage_r_3__result__63_, comp_stage_r_3__result__62_, comp_stage_r_3__result__61_, comp_stage_r_3__result__60_, comp_stage_r_3__result__59_, comp_stage_r_3__result__58_, comp_stage_r_3__result__57_, comp_stage_r_3__result__56_, comp_stage_r_3__result__55_, comp_stage_r_3__result__54_, comp_stage_r_3__result__53_, comp_stage_r_3__result__52_, comp_stage_r_3__result__51_, comp_stage_r_3__result__50_, comp_stage_r_3__result__49_, comp_stage_r_3__result__48_, comp_stage_r_3__result__47_, comp_stage_r_3__result__46_, comp_stage_r_3__result__45_, comp_stage_r_3__result__44_, comp_stage_r_3__result__43_, comp_stage_r_3__result__42_, comp_stage_r_3__result__41_, comp_stage_r_3__result__40_, comp_stage_r_3__result__39_, comp_stage_r_3__result__38_, comp_stage_r_3__result__37_, comp_stage_r_3__result__36_, comp_stage_r_3__result__35_, comp_stage_r_3__result__34_, comp_stage_r_3__result__33_, comp_stage_r_3__result__32_, comp_stage_r_3__result__31_, comp_stage_r_3__result__30_, comp_stage_r_3__result__29_, comp_stage_r_3__result__28_, comp_stage_r_3__result__27_, comp_stage_r_3__result__26_, comp_stage_r_3__result__25_, comp_stage_r_3__result__24_, comp_stage_r_3__result__23_, comp_stage_r_3__result__22_, comp_stage_r_3__result__21_, comp_stage_r_3__result__20_, comp_stage_r_3__result__19_, comp_stage_r_3__result__18_, comp_stage_r_3__result__17_, comp_stage_r_3__result__16_, comp_stage_r_3__result__15_, comp_stage_r_3__result__14_, comp_stage_r_3__result__13_, comp_stage_r_3__result__12_, comp_stage_r_3__result__11_, comp_stage_r_3__result__10_, comp_stage_r_3__result__9_, comp_stage_r_3__result__8_, comp_stage_r_3__result__7_, comp_stage_r_3__result__6_, comp_stage_r_3__result__5_, comp_stage_r_3__result__4_, comp_stage_r_3__result__3_, comp_stage_r_3__result__2_, comp_stage_r_3__result__1_, comp_stage_r_3__result__0_, comp_stage_r_3__br_tgt__63_, comp_stage_r_3__br_tgt__62_, comp_stage_r_3__br_tgt__61_, comp_stage_r_3__br_tgt__60_, comp_stage_r_3__br_tgt__59_, comp_stage_r_3__br_tgt__58_, comp_stage_r_3__br_tgt__57_, comp_stage_r_3__br_tgt__56_, comp_stage_r_3__br_tgt__55_, comp_stage_r_3__br_tgt__54_, comp_stage_r_3__br_tgt__53_, comp_stage_r_3__br_tgt__52_, comp_stage_r_3__br_tgt__51_, comp_stage_r_3__br_tgt__50_, comp_stage_r_3__br_tgt__49_, comp_stage_r_3__br_tgt__48_, comp_stage_r_3__br_tgt__47_, comp_stage_r_3__br_tgt__46_, comp_stage_r_3__br_tgt__45_, comp_stage_r_3__br_tgt__44_, comp_stage_r_3__br_tgt__43_, comp_stage_r_3__br_tgt__42_, comp_stage_r_3__br_tgt__41_, comp_stage_r_3__br_tgt__40_, comp_stage_r_3__br_tgt__39_, comp_stage_r_3__br_tgt__38_, comp_stage_r_3__br_tgt__37_, comp_stage_r_3__br_tgt__36_, comp_stage_r_3__br_tgt__35_, comp_stage_r_3__br_tgt__34_, comp_stage_r_3__br_tgt__33_, comp_stage_r_3__br_tgt__32_, comp_stage_r_3__br_tgt__31_, comp_stage_r_3__br_tgt__30_, comp_stage_r_3__br_tgt__29_, comp_stage_r_3__br_tgt__28_, comp_stage_r_3__br_tgt__27_, comp_stage_r_3__br_tgt__26_, comp_stage_r_3__br_tgt__25_, comp_stage_r_3__br_tgt__24_, comp_stage_r_3__br_tgt__23_, comp_stage_r_3__br_tgt__22_, comp_stage_r_3__br_tgt__21_, comp_stage_r_3__br_tgt__20_, comp_stage_r_3__br_tgt__19_, comp_stage_r_3__br_tgt__18_, comp_stage_r_3__br_tgt__17_, comp_stage_r_3__br_tgt__16_, comp_stage_r_3__br_tgt__15_, comp_stage_r_3__br_tgt__14_, comp_stage_r_3__br_tgt__13_, comp_stage_r_3__br_tgt__12_, comp_stage_r_3__br_tgt__11_, comp_stage_r_3__br_tgt__10_, comp_stage_r_3__br_tgt__9_, comp_stage_r_3__br_tgt__8_, comp_stage_r_3__br_tgt__7_, comp_stage_r_3__br_tgt__6_, comp_stage_r_3__br_tgt__5_, comp_stage_r_3__br_tgt__4_, comp_stage_r_3__br_tgt__3_, comp_stage_r_3__br_tgt__2_, comp_stage_r_3__br_tgt__1_, comp_stage_r_3__br_tgt__0_, comp_stage_r_2__result__63_, comp_stage_r_2__result__62_, comp_stage_r_2__result__61_, comp_stage_r_2__result__60_, comp_stage_r_2__result__59_, comp_stage_r_2__result__58_, comp_stage_r_2__result__57_, comp_stage_r_2__result__56_, comp_stage_r_2__result__55_, comp_stage_r_2__result__54_, comp_stage_r_2__result__53_, comp_stage_r_2__result__52_, comp_stage_r_2__result__51_, comp_stage_r_2__result__50_, comp_stage_r_2__result__49_, comp_stage_r_2__result__48_, comp_stage_r_2__result__47_, comp_stage_r_2__result__46_, comp_stage_r_2__result__45_, comp_stage_r_2__result__44_, comp_stage_r_2__result__43_, comp_stage_r_2__result__42_, comp_stage_r_2__result__41_, comp_stage_r_2__result__40_, comp_stage_r_2__result__39_, comp_stage_r_2__result__38_, comp_stage_r_2__result__37_, comp_stage_r_2__result__36_, comp_stage_r_2__result__35_, comp_stage_r_2__result__34_, comp_stage_r_2__result__33_, comp_stage_r_2__result__32_, comp_stage_r_2__result__31_, comp_stage_r_2__result__30_, comp_stage_r_2__result__29_, comp_stage_r_2__result__28_, comp_stage_r_2__result__27_, comp_stage_r_2__result__26_, comp_stage_r_2__result__25_, comp_stage_r_2__result__24_, comp_stage_r_2__result__23_, comp_stage_r_2__result__22_, comp_stage_r_2__result__21_, comp_stage_r_2__result__20_, comp_stage_r_2__result__19_, comp_stage_r_2__result__18_, comp_stage_r_2__result__17_, comp_stage_r_2__result__16_, comp_stage_r_2__result__15_, comp_stage_r_2__result__14_, comp_stage_r_2__result__13_, comp_stage_r_2__result__12_, comp_stage_r_2__result__11_, comp_stage_r_2__result__10_, comp_stage_r_2__result__9_, comp_stage_r_2__result__8_, comp_stage_r_2__result__7_, comp_stage_r_2__result__6_, comp_stage_r_2__result__5_, comp_stage_r_2__result__4_, comp_stage_r_2__result__3_, comp_stage_r_2__result__2_, comp_stage_r_2__result__1_, comp_stage_r_2__result__0_, comp_stage_r_2__br_tgt__63_, comp_stage_r_2__br_tgt__62_, comp_stage_r_2__br_tgt__61_, comp_stage_r_2__br_tgt__60_, comp_stage_r_2__br_tgt__59_, comp_stage_r_2__br_tgt__58_, comp_stage_r_2__br_tgt__57_, comp_stage_r_2__br_tgt__56_, comp_stage_r_2__br_tgt__55_, comp_stage_r_2__br_tgt__54_, comp_stage_r_2__br_tgt__53_, comp_stage_r_2__br_tgt__52_, comp_stage_r_2__br_tgt__51_, comp_stage_r_2__br_tgt__50_, comp_stage_r_2__br_tgt__49_, comp_stage_r_2__br_tgt__48_, comp_stage_r_2__br_tgt__47_, comp_stage_r_2__br_tgt__46_, comp_stage_r_2__br_tgt__45_, comp_stage_r_2__br_tgt__44_, comp_stage_r_2__br_tgt__43_, comp_stage_r_2__br_tgt__42_, comp_stage_r_2__br_tgt__41_, comp_stage_r_2__br_tgt__40_, comp_stage_r_2__br_tgt__39_, comp_stage_r_2__br_tgt__38_, comp_stage_r_2__br_tgt__37_, comp_stage_r_2__br_tgt__36_, comp_stage_r_2__br_tgt__35_, comp_stage_r_2__br_tgt__34_, comp_stage_r_2__br_tgt__33_, comp_stage_r_2__br_tgt__32_, comp_stage_r_2__br_tgt__31_, comp_stage_r_2__br_tgt__30_, comp_stage_r_2__br_tgt__29_, comp_stage_r_2__br_tgt__28_, comp_stage_r_2__br_tgt__27_, comp_stage_r_2__br_tgt__26_, comp_stage_r_2__br_tgt__25_, comp_stage_r_2__br_tgt__24_, comp_stage_r_2__br_tgt__23_, comp_stage_r_2__br_tgt__22_, comp_stage_r_2__br_tgt__21_, comp_stage_r_2__br_tgt__20_, comp_stage_r_2__br_tgt__19_, comp_stage_r_2__br_tgt__18_, comp_stage_r_2__br_tgt__17_, comp_stage_r_2__br_tgt__16_, comp_stage_r_2__br_tgt__15_, comp_stage_r_2__br_tgt__14_, comp_stage_r_2__br_tgt__13_, comp_stage_r_2__br_tgt__12_, comp_stage_r_2__br_tgt__11_, comp_stage_r_2__br_tgt__10_, comp_stage_r_2__br_tgt__9_, comp_stage_r_2__br_tgt__8_, comp_stage_r_2__br_tgt__7_, comp_stage_r_2__br_tgt__6_, comp_stage_r_2__br_tgt__5_, comp_stage_r_2__br_tgt__4_, comp_stage_r_2__br_tgt__3_, comp_stage_r_2__br_tgt__2_, comp_stage_r_2__br_tgt__1_, comp_stage_r_2__br_tgt__0_, comp_stage_r_1__result__63_, comp_stage_r_1__result__62_, comp_stage_r_1__result__61_, comp_stage_r_1__result__60_, comp_stage_r_1__result__59_, comp_stage_r_1__result__58_, comp_stage_r_1__result__57_, comp_stage_r_1__result__56_, comp_stage_r_1__result__55_, comp_stage_r_1__result__54_, comp_stage_r_1__result__53_, comp_stage_r_1__result__52_, comp_stage_r_1__result__51_, comp_stage_r_1__result__50_, comp_stage_r_1__result__49_, comp_stage_r_1__result__48_, comp_stage_r_1__result__47_, comp_stage_r_1__result__46_, comp_stage_r_1__result__45_, comp_stage_r_1__result__44_, comp_stage_r_1__result__43_, comp_stage_r_1__result__42_, comp_stage_r_1__result__41_, comp_stage_r_1__result__40_, comp_stage_r_1__result__39_, comp_stage_r_1__result__38_, comp_stage_r_1__result__37_, comp_stage_r_1__result__36_, comp_stage_r_1__result__35_, comp_stage_r_1__result__34_, comp_stage_r_1__result__33_, comp_stage_r_1__result__32_, comp_stage_r_1__result__31_, comp_stage_r_1__result__30_, comp_stage_r_1__result__29_, comp_stage_r_1__result__28_, comp_stage_r_1__result__27_, comp_stage_r_1__result__26_, comp_stage_r_1__result__25_, comp_stage_r_1__result__24_, comp_stage_r_1__result__23_, comp_stage_r_1__result__22_, comp_stage_r_1__result__21_, comp_stage_r_1__result__20_, comp_stage_r_1__result__19_, comp_stage_r_1__result__18_, comp_stage_r_1__result__17_, comp_stage_r_1__result__16_, comp_stage_r_1__result__15_, comp_stage_r_1__result__14_, comp_stage_r_1__result__13_, comp_stage_r_1__result__12_, comp_stage_r_1__result__11_, comp_stage_r_1__result__10_, comp_stage_r_1__result__9_, comp_stage_r_1__result__8_, comp_stage_r_1__result__7_, comp_stage_r_1__result__6_, comp_stage_r_1__result__5_, comp_stage_r_1__result__4_, comp_stage_r_1__result__3_, comp_stage_r_1__result__2_, comp_stage_r_1__result__1_, comp_stage_r_1__result__0_, comp_stage_r_1__br_tgt__63_, comp_stage_r_1__br_tgt__62_, comp_stage_r_1__br_tgt__61_, comp_stage_r_1__br_tgt__60_, comp_stage_r_1__br_tgt__59_, comp_stage_r_1__br_tgt__58_, comp_stage_r_1__br_tgt__57_, comp_stage_r_1__br_tgt__56_, comp_stage_r_1__br_tgt__55_, comp_stage_r_1__br_tgt__54_, comp_stage_r_1__br_tgt__53_, comp_stage_r_1__br_tgt__52_, comp_stage_r_1__br_tgt__51_, comp_stage_r_1__br_tgt__50_, comp_stage_r_1__br_tgt__49_, comp_stage_r_1__br_tgt__48_, comp_stage_r_1__br_tgt__47_, comp_stage_r_1__br_tgt__46_, comp_stage_r_1__br_tgt__45_, comp_stage_r_1__br_tgt__44_, comp_stage_r_1__br_tgt__43_, comp_stage_r_1__br_tgt__42_, comp_stage_r_1__br_tgt__41_, comp_stage_r_1__br_tgt__40_, comp_stage_r_1__br_tgt__39_, comp_stage_r_1__br_tgt__38_, comp_stage_r_1__br_tgt__37_, comp_stage_r_1__br_tgt__36_, comp_stage_r_1__br_tgt__35_, comp_stage_r_1__br_tgt__34_, comp_stage_r_1__br_tgt__33_, comp_stage_r_1__br_tgt__32_, comp_stage_r_1__br_tgt__31_, comp_stage_r_1__br_tgt__30_, comp_stage_r_1__br_tgt__29_, comp_stage_r_1__br_tgt__28_, comp_stage_r_1__br_tgt__27_, comp_stage_r_1__br_tgt__26_, comp_stage_r_1__br_tgt__25_, comp_stage_r_1__br_tgt__24_, comp_stage_r_1__br_tgt__23_, comp_stage_r_1__br_tgt__22_, comp_stage_r_1__br_tgt__21_, comp_stage_r_1__br_tgt__20_, comp_stage_r_1__br_tgt__19_, comp_stage_r_1__br_tgt__18_, comp_stage_r_1__br_tgt__17_, comp_stage_r_1__br_tgt__16_, comp_stage_r_1__br_tgt__15_, comp_stage_r_1__br_tgt__14_, comp_stage_r_1__br_tgt__13_, comp_stage_r_1__br_tgt__12_, comp_stage_r_1__br_tgt__11_, comp_stage_r_1__br_tgt__10_, comp_stage_r_1__br_tgt__9_, comp_stage_r_1__br_tgt__8_, comp_stage_r_1__br_tgt__7_, comp_stage_r_1__br_tgt__6_, comp_stage_r_1__br_tgt__5_, comp_stage_r_1__br_tgt__4_, comp_stage_r_1__br_tgt__3_, comp_stage_r_1__br_tgt__2_, comp_stage_r_1__br_tgt__1_, comp_stage_r_1__br_tgt__0_, comp_stage_r_0__result__63_, comp_stage_r_0__result__62_, comp_stage_r_0__result__61_, comp_stage_r_0__result__60_, comp_stage_r_0__result__59_, comp_stage_r_0__result__58_, comp_stage_r_0__result__57_, comp_stage_r_0__result__56_, comp_stage_r_0__result__55_, comp_stage_r_0__result__54_, comp_stage_r_0__result__53_, comp_stage_r_0__result__52_, comp_stage_r_0__result__51_, comp_stage_r_0__result__50_, comp_stage_r_0__result__49_, comp_stage_r_0__result__48_, comp_stage_r_0__result__47_, comp_stage_r_0__result__46_, comp_stage_r_0__result__45_, comp_stage_r_0__result__44_, comp_stage_r_0__result__43_, comp_stage_r_0__result__42_, comp_stage_r_0__result__41_, comp_stage_r_0__result__40_, comp_stage_r_0__result__39_, comp_stage_r_0__result__38_, comp_stage_r_0__result__37_, comp_stage_r_0__result__36_, comp_stage_r_0__result__35_, comp_stage_r_0__result__34_, comp_stage_r_0__result__33_, comp_stage_r_0__result__32_, comp_stage_r_0__result__31_, comp_stage_r_0__result__30_, comp_stage_r_0__result__29_, comp_stage_r_0__result__28_, comp_stage_r_0__result__27_, comp_stage_r_0__result__26_, comp_stage_r_0__result__25_, comp_stage_r_0__result__24_, comp_stage_r_0__result__23_, comp_stage_r_0__result__22_, comp_stage_r_0__result__21_, comp_stage_r_0__result__20_, comp_stage_r_0__result__19_, comp_stage_r_0__result__18_, comp_stage_r_0__result__17_, comp_stage_r_0__result__16_, comp_stage_r_0__result__15_, comp_stage_r_0__result__14_, comp_stage_r_0__result__13_, comp_stage_r_0__result__12_, comp_stage_r_0__result__11_, comp_stage_r_0__result__10_, comp_stage_r_0__result__9_, comp_stage_r_0__result__8_, comp_stage_r_0__result__7_, comp_stage_r_0__result__6_, comp_stage_r_0__result__5_, comp_stage_r_0__result__4_, comp_stage_r_0__result__3_, comp_stage_r_0__result__2_, comp_stage_r_0__result__1_, comp_stage_r_0__result__0_, comp_stage_r_0__br_tgt__63_, comp_stage_r_0__br_tgt__62_, comp_stage_r_0__br_tgt__61_, comp_stage_r_0__br_tgt__60_, comp_stage_r_0__br_tgt__59_, comp_stage_r_0__br_tgt__58_, comp_stage_r_0__br_tgt__57_, comp_stage_r_0__br_tgt__56_, comp_stage_r_0__br_tgt__55_, comp_stage_r_0__br_tgt__54_, comp_stage_r_0__br_tgt__53_, comp_stage_r_0__br_tgt__52_, comp_stage_r_0__br_tgt__51_, comp_stage_r_0__br_tgt__50_, comp_stage_r_0__br_tgt__49_, comp_stage_r_0__br_tgt__48_, comp_stage_r_0__br_tgt__47_, comp_stage_r_0__br_tgt__46_, comp_stage_r_0__br_tgt__45_, comp_stage_r_0__br_tgt__44_, comp_stage_r_0__br_tgt__43_, comp_stage_r_0__br_tgt__42_, comp_stage_r_0__br_tgt__41_, comp_stage_r_0__br_tgt__40_, comp_stage_r_0__br_tgt__39_, comp_stage_r_0__br_tgt__38_, comp_stage_r_0__br_tgt__37_, comp_stage_r_0__br_tgt__36_, comp_stage_r_0__br_tgt__35_, comp_stage_r_0__br_tgt__34_, comp_stage_r_0__br_tgt__33_, comp_stage_r_0__br_tgt__32_, comp_stage_r_0__br_tgt__31_, comp_stage_r_0__br_tgt__30_, comp_stage_r_0__br_tgt__29_, comp_stage_r_0__br_tgt__28_, comp_stage_r_0__br_tgt__27_, comp_stage_r_0__br_tgt__26_, comp_stage_r_0__br_tgt__25_, comp_stage_r_0__br_tgt__24_, comp_stage_r_0__br_tgt__23_, comp_stage_r_0__br_tgt__22_, comp_stage_r_0__br_tgt__21_, comp_stage_r_0__br_tgt__20_, comp_stage_r_0__br_tgt__19_, comp_stage_r_0__br_tgt__18_, comp_stage_r_0__br_tgt__17_, comp_stage_r_0__br_tgt__16_, comp_stage_r_0__br_tgt__15_, comp_stage_r_0__br_tgt__14_, comp_stage_r_0__br_tgt__13_, comp_stage_r_0__br_tgt__12_, comp_stage_r_0__br_tgt__11_, comp_stage_r_0__br_tgt__10_, comp_stage_r_0__br_tgt__9_, comp_stage_r_0__br_tgt__8_, comp_stage_r_0__br_tgt__7_, comp_stage_r_0__br_tgt__6_, comp_stage_r_0__br_tgt__5_, comp_stage_r_0__br_tgt__4_, comp_stage_r_0__br_tgt__3_, comp_stage_r_0__br_tgt__2_, comp_stage_r_0__br_tgt__1_, comp_stage_r_0__br_tgt__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .data1_i({ fp_calc_result, mem_calc_result, mul_calc_result, int_calc_result_result__63_, int_calc_result_result__62_, int_calc_result_result__61_, int_calc_result_result__60_, int_calc_result_result__59_, int_calc_result_result__58_, int_calc_result_result__57_, int_calc_result_result__56_, int_calc_result_result__55_, int_calc_result_result__54_, int_calc_result_result__53_, int_calc_result_result__52_, int_calc_result_result__51_, int_calc_result_result__50_, int_calc_result_result__49_, int_calc_result_result__48_, int_calc_result_result__47_, int_calc_result_result__46_, int_calc_result_result__45_, int_calc_result_result__44_, int_calc_result_result__43_, int_calc_result_result__42_, int_calc_result_result__41_, int_calc_result_result__40_, int_calc_result_result__39_, int_calc_result_result__38_, int_calc_result_result__37_, int_calc_result_result__36_, int_calc_result_result__35_, int_calc_result_result__34_, int_calc_result_result__33_, int_calc_result_result__32_, int_calc_result_result__31_, int_calc_result_result__30_, int_calc_result_result__29_, int_calc_result_result__28_, int_calc_result_result__27_, int_calc_result_result__26_, int_calc_result_result__25_, int_calc_result_result__24_, int_calc_result_result__23_, int_calc_result_result__22_, int_calc_result_result__21_, int_calc_result_result__20_, int_calc_result_result__19_, int_calc_result_result__18_, int_calc_result_result__17_, int_calc_result_result__16_, int_calc_result_result__15_, int_calc_result_result__14_, int_calc_result_result__13_, int_calc_result_result__12_, int_calc_result_result__11_, int_calc_result_result__10_, int_calc_result_result__9_, int_calc_result_result__8_, int_calc_result_result__7_, int_calc_result_result__6_, int_calc_result_result__5_, int_calc_result_result__4_, int_calc_result_result__3_, int_calc_result_result__2_, int_calc_result_result__1_, int_calc_result_result__0_, calc_status_o[221:158], nop_calc_result }),
    .sel_i({ calc_stage_r_3__decode__pipe_fp_v_, calc_stage_r_2__decode__pipe_mem_v_, calc_stage_r_1__decode__pipe_mul_v_, calc_stage_r_0__decode__pipe_int_v_, 1'b1 }),
    .data_o(comp_stage_n)
  );


  bsg_dff_width_p640
  comp_stage_reg
  (
    .clk_i(clk_i),
    .data_i(comp_stage_n),
    .data_o({ cmt_trace_result_o, comp_stage_r_3__result__63_, comp_stage_r_3__result__62_, comp_stage_r_3__result__61_, comp_stage_r_3__result__60_, comp_stage_r_3__result__59_, comp_stage_r_3__result__58_, comp_stage_r_3__result__57_, comp_stage_r_3__result__56_, comp_stage_r_3__result__55_, comp_stage_r_3__result__54_, comp_stage_r_3__result__53_, comp_stage_r_3__result__52_, comp_stage_r_3__result__51_, comp_stage_r_3__result__50_, comp_stage_r_3__result__49_, comp_stage_r_3__result__48_, comp_stage_r_3__result__47_, comp_stage_r_3__result__46_, comp_stage_r_3__result__45_, comp_stage_r_3__result__44_, comp_stage_r_3__result__43_, comp_stage_r_3__result__42_, comp_stage_r_3__result__41_, comp_stage_r_3__result__40_, comp_stage_r_3__result__39_, comp_stage_r_3__result__38_, comp_stage_r_3__result__37_, comp_stage_r_3__result__36_, comp_stage_r_3__result__35_, comp_stage_r_3__result__34_, comp_stage_r_3__result__33_, comp_stage_r_3__result__32_, comp_stage_r_3__result__31_, comp_stage_r_3__result__30_, comp_stage_r_3__result__29_, comp_stage_r_3__result__28_, comp_stage_r_3__result__27_, comp_stage_r_3__result__26_, comp_stage_r_3__result__25_, comp_stage_r_3__result__24_, comp_stage_r_3__result__23_, comp_stage_r_3__result__22_, comp_stage_r_3__result__21_, comp_stage_r_3__result__20_, comp_stage_r_3__result__19_, comp_stage_r_3__result__18_, comp_stage_r_3__result__17_, comp_stage_r_3__result__16_, comp_stage_r_3__result__15_, comp_stage_r_3__result__14_, comp_stage_r_3__result__13_, comp_stage_r_3__result__12_, comp_stage_r_3__result__11_, comp_stage_r_3__result__10_, comp_stage_r_3__result__9_, comp_stage_r_3__result__8_, comp_stage_r_3__result__7_, comp_stage_r_3__result__6_, comp_stage_r_3__result__5_, comp_stage_r_3__result__4_, comp_stage_r_3__result__3_, comp_stage_r_3__result__2_, comp_stage_r_3__result__1_, comp_stage_r_3__result__0_, comp_stage_r_3__br_tgt__63_, comp_stage_r_3__br_tgt__62_, comp_stage_r_3__br_tgt__61_, comp_stage_r_3__br_tgt__60_, comp_stage_r_3__br_tgt__59_, comp_stage_r_3__br_tgt__58_, comp_stage_r_3__br_tgt__57_, comp_stage_r_3__br_tgt__56_, comp_stage_r_3__br_tgt__55_, comp_stage_r_3__br_tgt__54_, comp_stage_r_3__br_tgt__53_, comp_stage_r_3__br_tgt__52_, comp_stage_r_3__br_tgt__51_, comp_stage_r_3__br_tgt__50_, comp_stage_r_3__br_tgt__49_, comp_stage_r_3__br_tgt__48_, comp_stage_r_3__br_tgt__47_, comp_stage_r_3__br_tgt__46_, comp_stage_r_3__br_tgt__45_, comp_stage_r_3__br_tgt__44_, comp_stage_r_3__br_tgt__43_, comp_stage_r_3__br_tgt__42_, comp_stage_r_3__br_tgt__41_, comp_stage_r_3__br_tgt__40_, comp_stage_r_3__br_tgt__39_, comp_stage_r_3__br_tgt__38_, comp_stage_r_3__br_tgt__37_, comp_stage_r_3__br_tgt__36_, comp_stage_r_3__br_tgt__35_, comp_stage_r_3__br_tgt__34_, comp_stage_r_3__br_tgt__33_, comp_stage_r_3__br_tgt__32_, comp_stage_r_3__br_tgt__31_, comp_stage_r_3__br_tgt__30_, comp_stage_r_3__br_tgt__29_, comp_stage_r_3__br_tgt__28_, comp_stage_r_3__br_tgt__27_, comp_stage_r_3__br_tgt__26_, comp_stage_r_3__br_tgt__25_, comp_stage_r_3__br_tgt__24_, comp_stage_r_3__br_tgt__23_, comp_stage_r_3__br_tgt__22_, comp_stage_r_3__br_tgt__21_, comp_stage_r_3__br_tgt__20_, comp_stage_r_3__br_tgt__19_, comp_stage_r_3__br_tgt__18_, comp_stage_r_3__br_tgt__17_, comp_stage_r_3__br_tgt__16_, comp_stage_r_3__br_tgt__15_, comp_stage_r_3__br_tgt__14_, comp_stage_r_3__br_tgt__13_, comp_stage_r_3__br_tgt__12_, comp_stage_r_3__br_tgt__11_, comp_stage_r_3__br_tgt__10_, comp_stage_r_3__br_tgt__9_, comp_stage_r_3__br_tgt__8_, comp_stage_r_3__br_tgt__7_, comp_stage_r_3__br_tgt__6_, comp_stage_r_3__br_tgt__5_, comp_stage_r_3__br_tgt__4_, comp_stage_r_3__br_tgt__3_, comp_stage_r_3__br_tgt__2_, comp_stage_r_3__br_tgt__1_, comp_stage_r_3__br_tgt__0_, comp_stage_r_2__result__63_, comp_stage_r_2__result__62_, comp_stage_r_2__result__61_, comp_stage_r_2__result__60_, comp_stage_r_2__result__59_, comp_stage_r_2__result__58_, comp_stage_r_2__result__57_, comp_stage_r_2__result__56_, comp_stage_r_2__result__55_, comp_stage_r_2__result__54_, comp_stage_r_2__result__53_, comp_stage_r_2__result__52_, comp_stage_r_2__result__51_, comp_stage_r_2__result__50_, comp_stage_r_2__result__49_, comp_stage_r_2__result__48_, comp_stage_r_2__result__47_, comp_stage_r_2__result__46_, comp_stage_r_2__result__45_, comp_stage_r_2__result__44_, comp_stage_r_2__result__43_, comp_stage_r_2__result__42_, comp_stage_r_2__result__41_, comp_stage_r_2__result__40_, comp_stage_r_2__result__39_, comp_stage_r_2__result__38_, comp_stage_r_2__result__37_, comp_stage_r_2__result__36_, comp_stage_r_2__result__35_, comp_stage_r_2__result__34_, comp_stage_r_2__result__33_, comp_stage_r_2__result__32_, comp_stage_r_2__result__31_, comp_stage_r_2__result__30_, comp_stage_r_2__result__29_, comp_stage_r_2__result__28_, comp_stage_r_2__result__27_, comp_stage_r_2__result__26_, comp_stage_r_2__result__25_, comp_stage_r_2__result__24_, comp_stage_r_2__result__23_, comp_stage_r_2__result__22_, comp_stage_r_2__result__21_, comp_stage_r_2__result__20_, comp_stage_r_2__result__19_, comp_stage_r_2__result__18_, comp_stage_r_2__result__17_, comp_stage_r_2__result__16_, comp_stage_r_2__result__15_, comp_stage_r_2__result__14_, comp_stage_r_2__result__13_, comp_stage_r_2__result__12_, comp_stage_r_2__result__11_, comp_stage_r_2__result__10_, comp_stage_r_2__result__9_, comp_stage_r_2__result__8_, comp_stage_r_2__result__7_, comp_stage_r_2__result__6_, comp_stage_r_2__result__5_, comp_stage_r_2__result__4_, comp_stage_r_2__result__3_, comp_stage_r_2__result__2_, comp_stage_r_2__result__1_, comp_stage_r_2__result__0_, comp_stage_r_2__br_tgt__63_, comp_stage_r_2__br_tgt__62_, comp_stage_r_2__br_tgt__61_, comp_stage_r_2__br_tgt__60_, comp_stage_r_2__br_tgt__59_, comp_stage_r_2__br_tgt__58_, comp_stage_r_2__br_tgt__57_, comp_stage_r_2__br_tgt__56_, comp_stage_r_2__br_tgt__55_, comp_stage_r_2__br_tgt__54_, comp_stage_r_2__br_tgt__53_, comp_stage_r_2__br_tgt__52_, comp_stage_r_2__br_tgt__51_, comp_stage_r_2__br_tgt__50_, comp_stage_r_2__br_tgt__49_, comp_stage_r_2__br_tgt__48_, comp_stage_r_2__br_tgt__47_, comp_stage_r_2__br_tgt__46_, comp_stage_r_2__br_tgt__45_, comp_stage_r_2__br_tgt__44_, comp_stage_r_2__br_tgt__43_, comp_stage_r_2__br_tgt__42_, comp_stage_r_2__br_tgt__41_, comp_stage_r_2__br_tgt__40_, comp_stage_r_2__br_tgt__39_, comp_stage_r_2__br_tgt__38_, comp_stage_r_2__br_tgt__37_, comp_stage_r_2__br_tgt__36_, comp_stage_r_2__br_tgt__35_, comp_stage_r_2__br_tgt__34_, comp_stage_r_2__br_tgt__33_, comp_stage_r_2__br_tgt__32_, comp_stage_r_2__br_tgt__31_, comp_stage_r_2__br_tgt__30_, comp_stage_r_2__br_tgt__29_, comp_stage_r_2__br_tgt__28_, comp_stage_r_2__br_tgt__27_, comp_stage_r_2__br_tgt__26_, comp_stage_r_2__br_tgt__25_, comp_stage_r_2__br_tgt__24_, comp_stage_r_2__br_tgt__23_, comp_stage_r_2__br_tgt__22_, comp_stage_r_2__br_tgt__21_, comp_stage_r_2__br_tgt__20_, comp_stage_r_2__br_tgt__19_, comp_stage_r_2__br_tgt__18_, comp_stage_r_2__br_tgt__17_, comp_stage_r_2__br_tgt__16_, comp_stage_r_2__br_tgt__15_, comp_stage_r_2__br_tgt__14_, comp_stage_r_2__br_tgt__13_, comp_stage_r_2__br_tgt__12_, comp_stage_r_2__br_tgt__11_, comp_stage_r_2__br_tgt__10_, comp_stage_r_2__br_tgt__9_, comp_stage_r_2__br_tgt__8_, comp_stage_r_2__br_tgt__7_, comp_stage_r_2__br_tgt__6_, comp_stage_r_2__br_tgt__5_, comp_stage_r_2__br_tgt__4_, comp_stage_r_2__br_tgt__3_, comp_stage_r_2__br_tgt__2_, comp_stage_r_2__br_tgt__1_, comp_stage_r_2__br_tgt__0_, comp_stage_r_1__result__63_, comp_stage_r_1__result__62_, comp_stage_r_1__result__61_, comp_stage_r_1__result__60_, comp_stage_r_1__result__59_, comp_stage_r_1__result__58_, comp_stage_r_1__result__57_, comp_stage_r_1__result__56_, comp_stage_r_1__result__55_, comp_stage_r_1__result__54_, comp_stage_r_1__result__53_, comp_stage_r_1__result__52_, comp_stage_r_1__result__51_, comp_stage_r_1__result__50_, comp_stage_r_1__result__49_, comp_stage_r_1__result__48_, comp_stage_r_1__result__47_, comp_stage_r_1__result__46_, comp_stage_r_1__result__45_, comp_stage_r_1__result__44_, comp_stage_r_1__result__43_, comp_stage_r_1__result__42_, comp_stage_r_1__result__41_, comp_stage_r_1__result__40_, comp_stage_r_1__result__39_, comp_stage_r_1__result__38_, comp_stage_r_1__result__37_, comp_stage_r_1__result__36_, comp_stage_r_1__result__35_, comp_stage_r_1__result__34_, comp_stage_r_1__result__33_, comp_stage_r_1__result__32_, comp_stage_r_1__result__31_, comp_stage_r_1__result__30_, comp_stage_r_1__result__29_, comp_stage_r_1__result__28_, comp_stage_r_1__result__27_, comp_stage_r_1__result__26_, comp_stage_r_1__result__25_, comp_stage_r_1__result__24_, comp_stage_r_1__result__23_, comp_stage_r_1__result__22_, comp_stage_r_1__result__21_, comp_stage_r_1__result__20_, comp_stage_r_1__result__19_, comp_stage_r_1__result__18_, comp_stage_r_1__result__17_, comp_stage_r_1__result__16_, comp_stage_r_1__result__15_, comp_stage_r_1__result__14_, comp_stage_r_1__result__13_, comp_stage_r_1__result__12_, comp_stage_r_1__result__11_, comp_stage_r_1__result__10_, comp_stage_r_1__result__9_, comp_stage_r_1__result__8_, comp_stage_r_1__result__7_, comp_stage_r_1__result__6_, comp_stage_r_1__result__5_, comp_stage_r_1__result__4_, comp_stage_r_1__result__3_, comp_stage_r_1__result__2_, comp_stage_r_1__result__1_, comp_stage_r_1__result__0_, comp_stage_r_1__br_tgt__63_, comp_stage_r_1__br_tgt__62_, comp_stage_r_1__br_tgt__61_, comp_stage_r_1__br_tgt__60_, comp_stage_r_1__br_tgt__59_, comp_stage_r_1__br_tgt__58_, comp_stage_r_1__br_tgt__57_, comp_stage_r_1__br_tgt__56_, comp_stage_r_1__br_tgt__55_, comp_stage_r_1__br_tgt__54_, comp_stage_r_1__br_tgt__53_, comp_stage_r_1__br_tgt__52_, comp_stage_r_1__br_tgt__51_, comp_stage_r_1__br_tgt__50_, comp_stage_r_1__br_tgt__49_, comp_stage_r_1__br_tgt__48_, comp_stage_r_1__br_tgt__47_, comp_stage_r_1__br_tgt__46_, comp_stage_r_1__br_tgt__45_, comp_stage_r_1__br_tgt__44_, comp_stage_r_1__br_tgt__43_, comp_stage_r_1__br_tgt__42_, comp_stage_r_1__br_tgt__41_, comp_stage_r_1__br_tgt__40_, comp_stage_r_1__br_tgt__39_, comp_stage_r_1__br_tgt__38_, comp_stage_r_1__br_tgt__37_, comp_stage_r_1__br_tgt__36_, comp_stage_r_1__br_tgt__35_, comp_stage_r_1__br_tgt__34_, comp_stage_r_1__br_tgt__33_, comp_stage_r_1__br_tgt__32_, comp_stage_r_1__br_tgt__31_, comp_stage_r_1__br_tgt__30_, comp_stage_r_1__br_tgt__29_, comp_stage_r_1__br_tgt__28_, comp_stage_r_1__br_tgt__27_, comp_stage_r_1__br_tgt__26_, comp_stage_r_1__br_tgt__25_, comp_stage_r_1__br_tgt__24_, comp_stage_r_1__br_tgt__23_, comp_stage_r_1__br_tgt__22_, comp_stage_r_1__br_tgt__21_, comp_stage_r_1__br_tgt__20_, comp_stage_r_1__br_tgt__19_, comp_stage_r_1__br_tgt__18_, comp_stage_r_1__br_tgt__17_, comp_stage_r_1__br_tgt__16_, comp_stage_r_1__br_tgt__15_, comp_stage_r_1__br_tgt__14_, comp_stage_r_1__br_tgt__13_, comp_stage_r_1__br_tgt__12_, comp_stage_r_1__br_tgt__11_, comp_stage_r_1__br_tgt__10_, comp_stage_r_1__br_tgt__9_, comp_stage_r_1__br_tgt__8_, comp_stage_r_1__br_tgt__7_, comp_stage_r_1__br_tgt__6_, comp_stage_r_1__br_tgt__5_, comp_stage_r_1__br_tgt__4_, comp_stage_r_1__br_tgt__3_, comp_stage_r_1__br_tgt__2_, comp_stage_r_1__br_tgt__1_, comp_stage_r_1__br_tgt__0_, comp_stage_r_0__result__63_, comp_stage_r_0__result__62_, comp_stage_r_0__result__61_, comp_stage_r_0__result__60_, comp_stage_r_0__result__59_, comp_stage_r_0__result__58_, comp_stage_r_0__result__57_, comp_stage_r_0__result__56_, comp_stage_r_0__result__55_, comp_stage_r_0__result__54_, comp_stage_r_0__result__53_, comp_stage_r_0__result__52_, comp_stage_r_0__result__51_, comp_stage_r_0__result__50_, comp_stage_r_0__result__49_, comp_stage_r_0__result__48_, comp_stage_r_0__result__47_, comp_stage_r_0__result__46_, comp_stage_r_0__result__45_, comp_stage_r_0__result__44_, comp_stage_r_0__result__43_, comp_stage_r_0__result__42_, comp_stage_r_0__result__41_, comp_stage_r_0__result__40_, comp_stage_r_0__result__39_, comp_stage_r_0__result__38_, comp_stage_r_0__result__37_, comp_stage_r_0__result__36_, comp_stage_r_0__result__35_, comp_stage_r_0__result__34_, comp_stage_r_0__result__33_, comp_stage_r_0__result__32_, comp_stage_r_0__result__31_, comp_stage_r_0__result__30_, comp_stage_r_0__result__29_, comp_stage_r_0__result__28_, comp_stage_r_0__result__27_, comp_stage_r_0__result__26_, comp_stage_r_0__result__25_, comp_stage_r_0__result__24_, comp_stage_r_0__result__23_, comp_stage_r_0__result__22_, comp_stage_r_0__result__21_, comp_stage_r_0__result__20_, comp_stage_r_0__result__19_, comp_stage_r_0__result__18_, comp_stage_r_0__result__17_, comp_stage_r_0__result__16_, comp_stage_r_0__result__15_, comp_stage_r_0__result__14_, comp_stage_r_0__result__13_, comp_stage_r_0__result__12_, comp_stage_r_0__result__11_, comp_stage_r_0__result__10_, comp_stage_r_0__result__9_, comp_stage_r_0__result__8_, comp_stage_r_0__result__7_, comp_stage_r_0__result__6_, comp_stage_r_0__result__5_, comp_stage_r_0__result__4_, comp_stage_r_0__result__3_, comp_stage_r_0__result__2_, comp_stage_r_0__result__1_, comp_stage_r_0__result__0_, comp_stage_r_0__br_tgt__63_, comp_stage_r_0__br_tgt__62_, comp_stage_r_0__br_tgt__61_, comp_stage_r_0__br_tgt__60_, comp_stage_r_0__br_tgt__59_, comp_stage_r_0__br_tgt__58_, comp_stage_r_0__br_tgt__57_, comp_stage_r_0__br_tgt__56_, comp_stage_r_0__br_tgt__55_, comp_stage_r_0__br_tgt__54_, comp_stage_r_0__br_tgt__53_, comp_stage_r_0__br_tgt__52_, comp_stage_r_0__br_tgt__51_, comp_stage_r_0__br_tgt__50_, comp_stage_r_0__br_tgt__49_, comp_stage_r_0__br_tgt__48_, comp_stage_r_0__br_tgt__47_, comp_stage_r_0__br_tgt__46_, comp_stage_r_0__br_tgt__45_, comp_stage_r_0__br_tgt__44_, comp_stage_r_0__br_tgt__43_, comp_stage_r_0__br_tgt__42_, comp_stage_r_0__br_tgt__41_, comp_stage_r_0__br_tgt__40_, comp_stage_r_0__br_tgt__39_, comp_stage_r_0__br_tgt__38_, comp_stage_r_0__br_tgt__37_, comp_stage_r_0__br_tgt__36_, comp_stage_r_0__br_tgt__35_, comp_stage_r_0__br_tgt__34_, comp_stage_r_0__br_tgt__33_, comp_stage_r_0__br_tgt__32_, comp_stage_r_0__br_tgt__31_, comp_stage_r_0__br_tgt__30_, comp_stage_r_0__br_tgt__29_, comp_stage_r_0__br_tgt__28_, comp_stage_r_0__br_tgt__27_, comp_stage_r_0__br_tgt__26_, comp_stage_r_0__br_tgt__25_, comp_stage_r_0__br_tgt__24_, comp_stage_r_0__br_tgt__23_, comp_stage_r_0__br_tgt__22_, comp_stage_r_0__br_tgt__21_, comp_stage_r_0__br_tgt__20_, comp_stage_r_0__br_tgt__19_, comp_stage_r_0__br_tgt__18_, comp_stage_r_0__br_tgt__17_, comp_stage_r_0__br_tgt__16_, comp_stage_r_0__br_tgt__15_, comp_stage_r_0__br_tgt__14_, comp_stage_r_0__br_tgt__13_, comp_stage_r_0__br_tgt__12_, comp_stage_r_0__br_tgt__11_, comp_stage_r_0__br_tgt__10_, comp_stage_r_0__br_tgt__9_, comp_stage_r_0__br_tgt__8_, comp_stage_r_0__br_tgt__7_, comp_stage_r_0__br_tgt__6_, comp_stage_r_0__br_tgt__5_, comp_stage_r_0__br_tgt__4_, comp_stage_r_0__br_tgt__3_, comp_stage_r_0__br_tgt__2_, comp_stage_r_0__br_tgt__1_, comp_stage_r_0__br_tgt__0_ })
  );


  bsg_dff_width_p35
  exc_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ exc_stage_r_3__poison_v_, exc_stage_r_3__roll_v_, exc_stage_r_3__illegal_instr_v_, exc_stage_r_3__tlb_miss_v_, exc_stage_r_3__load_fault_v_, exc_stage_r_3__store_fault_v_, exc_stage_r_3__cache_miss_v_, exc_stage_r_2__poison_v_, exc_stage_n_3__roll_v_, exc_stage_r_2__illegal_instr_v_, exc_stage_r_2__tlb_miss_v_, exc_stage_r_2__load_fault_v_, exc_stage_r_2__store_fault_v_, exc_stage_n_3__cache_miss_v_, exc_stage_n_2__poison_v_, exc_stage_n_2__roll_v_, exc_stage_r_1__illegal_instr_v_, exc_stage_r_1__tlb_miss_v_, exc_stage_r_1__load_fault_v_, exc_stage_r_1__store_fault_v_, exc_stage_r_1__cache_miss_v_, exc_stage_n_1__poison_v_, exc_stage_n_1__roll_v_, exc_stage_r_0__illegal_instr_v_, exc_stage_r_0__tlb_miss_v_, exc_stage_r_0__load_fault_v_, exc_stage_r_0__store_fault_v_, exc_stage_r_0__cache_miss_v_, chk_poison_isd_i, chk_roll_i, exc_stage_n_0__illegal_instr_v_, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .data_o({ cmt_trace_exc_o, exc_stage_r_3__poison_v_, exc_stage_r_3__roll_v_, exc_stage_r_3__illegal_instr_v_, exc_stage_r_3__tlb_miss_v_, exc_stage_r_3__load_fault_v_, exc_stage_r_3__store_fault_v_, exc_stage_r_3__cache_miss_v_, exc_stage_r_2__poison_v_, exc_stage_r_2__roll_v_, exc_stage_r_2__illegal_instr_v_, exc_stage_r_2__tlb_miss_v_, exc_stage_r_2__load_fault_v_, exc_stage_r_2__store_fault_v_, exc_stage_r_2__cache_miss_v_, exc_stage_r_1__poison_v_, exc_stage_r_1__roll_v_, exc_stage_r_1__illegal_instr_v_, exc_stage_r_1__tlb_miss_v_, exc_stage_r_1__load_fault_v_, exc_stage_r_1__store_fault_v_, exc_stage_r_1__cache_miss_v_, exc_stage_r_0__poison_v_, exc_stage_r_0__roll_v_, exc_stage_r_0__illegal_instr_v_, exc_stage_r_0__tlb_miss_v_, exc_stage_r_0__load_fault_v_, exc_stage_r_0__store_fault_v_, exc_stage_r_0__cache_miss_v_ })
  );

  assign issue_pkt_ready_o = N3 & N4;
  assign N3 = N1 & N2;
  assign N1 = chk_dispatch_v_i | N0;
  assign N0 = ~calc_status_o[301];
  assign N2 = ~chk_roll_i;
  assign N4 = ~chk_poison_isd_i;
  assign n_0_net_ = calc_stage_r_3__decode__irf_w_v_ & N11;
  assign N11 = ~N10;
  assign N10 = N9 | exc_stage_r_3__cache_miss_v_;
  assign N9 = N8 | exc_stage_r_3__store_fault_v_;
  assign N8 = N7 | exc_stage_r_3__load_fault_v_;
  assign N7 = N6 | exc_stage_r_3__tlb_miss_v_;
  assign N6 = N5 | exc_stage_r_3__illegal_instr_v_;
  assign N5 = exc_stage_r_3__poison_v_ | exc_stage_r_3__roll_v_;
  assign n_7_net_ = cmt_trace_stage_reg_o[32] & N18;
  assign N18 = ~N17;
  assign N17 = N16 | cmt_trace_exc_o[0];
  assign N16 = N15 | cmt_trace_exc_o[1];
  assign N15 = N14 | cmt_trace_exc_o[2];
  assign N14 = N13 | cmt_trace_exc_o[3];
  assign N13 = N12 | cmt_trace_exc_o[4];
  assign N12 = cmt_trace_exc_o[6] | cmt_trace_exc_o[5];
  assign n_15_net_ = issue_pkt_v_i | chk_dispatch_v_i;
  assign n_14_net_ = reset_i | chk_roll_i;
  assign n_17_net_ = issue_pkt_v_i | chk_dispatch_v_i;
  assign n_16_net_ = reset_i | chk_roll_i;
  assign n_20_net_ = N19 & N20;
  assign N19 = ~chk_dispatch_v_i;
  assign N20 = ~mmu_cmd_ready_i;
  assign n_19_net_ = N21 & mmu_cmd_ready_i;
  assign N21 = ~chk_dispatch_v_i;
  assign n_18_net_ = ~calc_status_o[301];
  assign calc_status_o[222] = calc_stage_r_0__decode__pipe_int_v_ & N28;
  assign N28 = ~N27;
  assign N27 = N26 | exc_stage_r_0__cache_miss_v_;
  assign N26 = N25 | exc_stage_r_0__store_fault_v_;
  assign N25 = N24 | exc_stage_r_0__load_fault_v_;
  assign N24 = N23 | exc_stage_r_0__tlb_miss_v_;
  assign N23 = N22 | exc_stage_r_0__illegal_instr_v_;
  assign N22 = exc_stage_r_0__poison_v_ | exc_stage_r_0__roll_v_;
  assign calc_status_o[120] = N29 | calc_stage_r_0__decode__jmp_v_;
  assign N29 = calc_stage_r_0__decode__br_v_ & int_calc_result_result__0_;
  assign calc_status_o[121] = calc_stage_r_0__decode__br_v_ | calc_stage_r_0__decode__jmp_v_;
  assign calc_status_o[119] = calc_stage_r_0__decode__instr_v_ & N36;
  assign N36 = ~N35;
  assign N35 = N34 | exc_stage_r_0__cache_miss_v_;
  assign N34 = N33 | exc_stage_r_0__store_fault_v_;
  assign N33 = N32 | exc_stage_r_0__load_fault_v_;
  assign N32 = N31 | exc_stage_r_0__tlb_miss_v_;
  assign N31 = N30 | exc_stage_r_0__illegal_instr_v_;
  assign N30 = exc_stage_r_0__poison_v_ | exc_stage_r_0__roll_v_;
  assign calc_status_o[78] = N44 & calc_stage_r_0__decode__irf_w_v_;
  assign N44 = calc_stage_r_0__decode__pipe_int_v_ & N43;
  assign N43 = ~N42;
  assign N42 = N41 | exc_stage_r_0__cache_miss_v_;
  assign N41 = N40 | exc_stage_r_0__store_fault_v_;
  assign N40 = N39 | exc_stage_r_0__load_fault_v_;
  assign N39 = N38 | exc_stage_r_0__tlb_miss_v_;
  assign N38 = N37 | exc_stage_r_0__illegal_instr_v_;
  assign N37 = exc_stage_r_0__poison_v_ | exc_stage_r_0__roll_v_;
  assign calc_status_o[77] = N52 & calc_stage_r_0__decode__irf_w_v_;
  assign N52 = calc_stage_r_0__decode__pipe_mul_v_ & N51;
  assign N51 = ~N50;
  assign N50 = N49 | exc_stage_r_0__cache_miss_v_;
  assign N49 = N48 | exc_stage_r_0__store_fault_v_;
  assign N48 = N47 | exc_stage_r_0__load_fault_v_;
  assign N47 = N46 | exc_stage_r_0__tlb_miss_v_;
  assign N46 = N45 | exc_stage_r_0__illegal_instr_v_;
  assign N45 = exc_stage_r_0__poison_v_ | exc_stage_r_0__roll_v_;
  assign calc_status_o[76] = N60 & calc_stage_r_0__decode__irf_w_v_;
  assign N60 = calc_stage_r_0__decode__pipe_mem_v_ & N59;
  assign N59 = ~N58;
  assign N58 = N57 | exc_stage_r_0__cache_miss_v_;
  assign N57 = N56 | exc_stage_r_0__store_fault_v_;
  assign N56 = N55 | exc_stage_r_0__load_fault_v_;
  assign N55 = N54 | exc_stage_r_0__tlb_miss_v_;
  assign N54 = N53 | exc_stage_r_0__illegal_instr_v_;
  assign N53 = exc_stage_r_0__poison_v_ | exc_stage_r_0__roll_v_;
  assign calc_status_o[75] = N68 & calc_stage_r_0__decode__frf_w_v_;
  assign N68 = calc_stage_r_0__decode__pipe_mem_v_ & N67;
  assign N67 = ~N66;
  assign N66 = N65 | exc_stage_r_0__cache_miss_v_;
  assign N65 = N64 | exc_stage_r_0__store_fault_v_;
  assign N64 = N63 | exc_stage_r_0__load_fault_v_;
  assign N63 = N62 | exc_stage_r_0__tlb_miss_v_;
  assign N62 = N61 | exc_stage_r_0__illegal_instr_v_;
  assign N61 = exc_stage_r_0__poison_v_ | exc_stage_r_0__roll_v_;
  assign calc_status_o[74] = N76 & calc_stage_r_0__decode__frf_w_v_;
  assign N76 = calc_stage_r_0__decode__pipe_fp_v_ & N75;
  assign N75 = ~N74;
  assign N74 = N73 | exc_stage_r_0__cache_miss_v_;
  assign N73 = N72 | exc_stage_r_0__store_fault_v_;
  assign N72 = N71 | exc_stage_r_0__load_fault_v_;
  assign N71 = N70 | exc_stage_r_0__tlb_miss_v_;
  assign N70 = N69 | exc_stage_r_0__illegal_instr_v_;
  assign N69 = exc_stage_r_0__poison_v_ | exc_stage_r_0__roll_v_;
  assign calc_status_o[88] = N84 & calc_stage_r_1__decode__irf_w_v_;
  assign N84 = calc_stage_r_1__decode__pipe_int_v_ & N83;
  assign N83 = ~N82;
  assign N82 = N81 | exc_stage_r_1__cache_miss_v_;
  assign N81 = N80 | exc_stage_r_1__store_fault_v_;
  assign N80 = N79 | exc_stage_r_1__load_fault_v_;
  assign N79 = N78 | exc_stage_r_1__tlb_miss_v_;
  assign N78 = N77 | exc_stage_r_1__illegal_instr_v_;
  assign N77 = exc_stage_r_1__poison_v_ | exc_stage_r_1__roll_v_;
  assign calc_status_o[87] = N92 & calc_stage_r_1__decode__irf_w_v_;
  assign N92 = calc_stage_r_1__decode__pipe_mul_v_ & N91;
  assign N91 = ~N90;
  assign N90 = N89 | exc_stage_r_1__cache_miss_v_;
  assign N89 = N88 | exc_stage_r_1__store_fault_v_;
  assign N88 = N87 | exc_stage_r_1__load_fault_v_;
  assign N87 = N86 | exc_stage_r_1__tlb_miss_v_;
  assign N86 = N85 | exc_stage_r_1__illegal_instr_v_;
  assign N85 = exc_stage_r_1__poison_v_ | exc_stage_r_1__roll_v_;
  assign calc_status_o[86] = N100 & calc_stage_r_1__decode__irf_w_v_;
  assign N100 = calc_stage_r_1__decode__pipe_mem_v_ & N99;
  assign N99 = ~N98;
  assign N98 = N97 | exc_stage_r_1__cache_miss_v_;
  assign N97 = N96 | exc_stage_r_1__store_fault_v_;
  assign N96 = N95 | exc_stage_r_1__load_fault_v_;
  assign N95 = N94 | exc_stage_r_1__tlb_miss_v_;
  assign N94 = N93 | exc_stage_r_1__illegal_instr_v_;
  assign N93 = exc_stage_r_1__poison_v_ | exc_stage_r_1__roll_v_;
  assign calc_status_o[85] = N108 & calc_stage_r_1__decode__frf_w_v_;
  assign N108 = calc_stage_r_1__decode__pipe_mem_v_ & N107;
  assign N107 = ~N106;
  assign N106 = N105 | exc_stage_r_1__cache_miss_v_;
  assign N105 = N104 | exc_stage_r_1__store_fault_v_;
  assign N104 = N103 | exc_stage_r_1__load_fault_v_;
  assign N103 = N102 | exc_stage_r_1__tlb_miss_v_;
  assign N102 = N101 | exc_stage_r_1__illegal_instr_v_;
  assign N101 = exc_stage_r_1__poison_v_ | exc_stage_r_1__roll_v_;
  assign calc_status_o[84] = N116 & calc_stage_r_1__decode__frf_w_v_;
  assign N116 = calc_stage_r_1__decode__pipe_fp_v_ & N115;
  assign N115 = ~N114;
  assign N114 = N113 | exc_stage_r_1__cache_miss_v_;
  assign N113 = N112 | exc_stage_r_1__store_fault_v_;
  assign N112 = N111 | exc_stage_r_1__load_fault_v_;
  assign N111 = N110 | exc_stage_r_1__tlb_miss_v_;
  assign N110 = N109 | exc_stage_r_1__illegal_instr_v_;
  assign N109 = exc_stage_r_1__poison_v_ | exc_stage_r_1__roll_v_;
  assign calc_status_o[98] = N124 & calc_stage_r_2__decode__irf_w_v_;
  assign N124 = calc_stage_r_2__decode__pipe_int_v_ & N123;
  assign N123 = ~N122;
  assign N122 = N121 | exc_stage_r_2__cache_miss_v_;
  assign N121 = N120 | exc_stage_r_2__store_fault_v_;
  assign N120 = N119 | exc_stage_r_2__load_fault_v_;
  assign N119 = N118 | exc_stage_r_2__tlb_miss_v_;
  assign N118 = N117 | exc_stage_r_2__illegal_instr_v_;
  assign N117 = exc_stage_r_2__poison_v_ | exc_stage_r_2__roll_v_;
  assign calc_status_o[97] = N132 & calc_stage_r_2__decode__irf_w_v_;
  assign N132 = calc_stage_r_2__decode__pipe_mul_v_ & N131;
  assign N131 = ~N130;
  assign N130 = N129 | exc_stage_r_2__cache_miss_v_;
  assign N129 = N128 | exc_stage_r_2__store_fault_v_;
  assign N128 = N127 | exc_stage_r_2__load_fault_v_;
  assign N127 = N126 | exc_stage_r_2__tlb_miss_v_;
  assign N126 = N125 | exc_stage_r_2__illegal_instr_v_;
  assign N125 = exc_stage_r_2__poison_v_ | exc_stage_r_2__roll_v_;
  assign calc_status_o[96] = N140 & calc_stage_r_2__decode__irf_w_v_;
  assign N140 = calc_stage_r_2__decode__pipe_mem_v_ & N139;
  assign N139 = ~N138;
  assign N138 = N137 | exc_stage_r_2__cache_miss_v_;
  assign N137 = N136 | exc_stage_r_2__store_fault_v_;
  assign N136 = N135 | exc_stage_r_2__load_fault_v_;
  assign N135 = N134 | exc_stage_r_2__tlb_miss_v_;
  assign N134 = N133 | exc_stage_r_2__illegal_instr_v_;
  assign N133 = exc_stage_r_2__poison_v_ | exc_stage_r_2__roll_v_;
  assign calc_status_o[95] = N148 & calc_stage_r_2__decode__frf_w_v_;
  assign N148 = calc_stage_r_2__decode__pipe_mem_v_ & N147;
  assign N147 = ~N146;
  assign N146 = N145 | exc_stage_r_2__cache_miss_v_;
  assign N145 = N144 | exc_stage_r_2__store_fault_v_;
  assign N144 = N143 | exc_stage_r_2__load_fault_v_;
  assign N143 = N142 | exc_stage_r_2__tlb_miss_v_;
  assign N142 = N141 | exc_stage_r_2__illegal_instr_v_;
  assign N141 = exc_stage_r_2__poison_v_ | exc_stage_r_2__roll_v_;
  assign calc_status_o[94] = N156 & calc_stage_r_2__decode__frf_w_v_;
  assign N156 = calc_stage_r_2__decode__pipe_fp_v_ & N155;
  assign N155 = ~N154;
  assign N154 = N153 | exc_stage_r_2__cache_miss_v_;
  assign N153 = N152 | exc_stage_r_2__store_fault_v_;
  assign N152 = N151 | exc_stage_r_2__load_fault_v_;
  assign N151 = N150 | exc_stage_r_2__tlb_miss_v_;
  assign N150 = N149 | exc_stage_r_2__illegal_instr_v_;
  assign N149 = exc_stage_r_2__poison_v_ | exc_stage_r_2__roll_v_;
  assign calc_status_o[108] = N164 & calc_stage_r_3__decode__irf_w_v_;
  assign N164 = calc_stage_r_3__decode__pipe_int_v_ & N163;
  assign N163 = ~N162;
  assign N162 = N161 | exc_stage_r_3__cache_miss_v_;
  assign N161 = N160 | exc_stage_r_3__store_fault_v_;
  assign N160 = N159 | exc_stage_r_3__load_fault_v_;
  assign N159 = N158 | exc_stage_r_3__tlb_miss_v_;
  assign N158 = N157 | exc_stage_r_3__illegal_instr_v_;
  assign N157 = exc_stage_r_3__poison_v_ | exc_stage_r_3__roll_v_;
  assign calc_status_o[107] = N172 & calc_stage_r_3__decode__irf_w_v_;
  assign N172 = calc_stage_r_3__decode__pipe_mul_v_ & N171;
  assign N171 = ~N170;
  assign N170 = N169 | exc_stage_r_3__cache_miss_v_;
  assign N169 = N168 | exc_stage_r_3__store_fault_v_;
  assign N168 = N167 | exc_stage_r_3__load_fault_v_;
  assign N167 = N166 | exc_stage_r_3__tlb_miss_v_;
  assign N166 = N165 | exc_stage_r_3__illegal_instr_v_;
  assign N165 = exc_stage_r_3__poison_v_ | exc_stage_r_3__roll_v_;
  assign calc_status_o[106] = N180 & calc_stage_r_3__decode__irf_w_v_;
  assign N180 = calc_stage_r_3__decode__pipe_mem_v_ & N179;
  assign N179 = ~N178;
  assign N178 = N177 | exc_stage_r_3__cache_miss_v_;
  assign N177 = N176 | exc_stage_r_3__store_fault_v_;
  assign N176 = N175 | exc_stage_r_3__load_fault_v_;
  assign N175 = N174 | exc_stage_r_3__tlb_miss_v_;
  assign N174 = N173 | exc_stage_r_3__illegal_instr_v_;
  assign N173 = exc_stage_r_3__poison_v_ | exc_stage_r_3__roll_v_;
  assign calc_status_o[105] = N188 & calc_stage_r_3__decode__frf_w_v_;
  assign N188 = calc_stage_r_3__decode__pipe_mem_v_ & N187;
  assign N187 = ~N186;
  assign N186 = N185 | exc_stage_r_3__cache_miss_v_;
  assign N185 = N184 | exc_stage_r_3__store_fault_v_;
  assign N184 = N183 | exc_stage_r_3__load_fault_v_;
  assign N183 = N182 | exc_stage_r_3__tlb_miss_v_;
  assign N182 = N181 | exc_stage_r_3__illegal_instr_v_;
  assign N181 = exc_stage_r_3__poison_v_ | exc_stage_r_3__roll_v_;
  assign calc_status_o[104] = N196 & calc_stage_r_3__decode__frf_w_v_;
  assign N196 = calc_stage_r_3__decode__pipe_fp_v_ & N195;
  assign N195 = ~N194;
  assign N194 = N193 | exc_stage_r_3__cache_miss_v_;
  assign N193 = N192 | exc_stage_r_3__store_fault_v_;
  assign N192 = N191 | exc_stage_r_3__load_fault_v_;
  assign N191 = N190 | exc_stage_r_3__tlb_miss_v_;
  assign N190 = N189 | exc_stage_r_3__illegal_instr_v_;
  assign N189 = exc_stage_r_3__poison_v_ | exc_stage_r_3__roll_v_;
  assign calc_status_o[118] = N204 & cmt_trace_stage_reg_o[33];
  assign N204 = cmt_trace_stage_reg_o[37] & N203;
  assign N203 = ~N202;
  assign N202 = N201 | cmt_trace_exc_o[0];
  assign N201 = N200 | cmt_trace_exc_o[1];
  assign N200 = N199 | cmt_trace_exc_o[2];
  assign N199 = N198 | cmt_trace_exc_o[3];
  assign N198 = N197 | cmt_trace_exc_o[4];
  assign N197 = cmt_trace_exc_o[6] | cmt_trace_exc_o[5];
  assign calc_status_o[117] = N212 & cmt_trace_stage_reg_o[33];
  assign N212 = cmt_trace_stage_reg_o[36] & N211;
  assign N211 = ~N210;
  assign N210 = N209 | cmt_trace_exc_o[0];
  assign N209 = N208 | cmt_trace_exc_o[1];
  assign N208 = N207 | cmt_trace_exc_o[2];
  assign N207 = N206 | cmt_trace_exc_o[3];
  assign N206 = N205 | cmt_trace_exc_o[4];
  assign N205 = cmt_trace_exc_o[6] | cmt_trace_exc_o[5];
  assign calc_status_o[116] = N220 & cmt_trace_stage_reg_o[33];
  assign N220 = cmt_trace_stage_reg_o[35] & N219;
  assign N219 = ~N218;
  assign N218 = N217 | cmt_trace_exc_o[0];
  assign N217 = N216 | cmt_trace_exc_o[1];
  assign N216 = N215 | cmt_trace_exc_o[2];
  assign N215 = N214 | cmt_trace_exc_o[3];
  assign N214 = N213 | cmt_trace_exc_o[4];
  assign N213 = cmt_trace_exc_o[6] | cmt_trace_exc_o[5];
  assign calc_status_o[115] = N228 & cmt_trace_stage_reg_o[32];
  assign N228 = cmt_trace_stage_reg_o[35] & N227;
  assign N227 = ~N226;
  assign N226 = N225 | cmt_trace_exc_o[0];
  assign N225 = N224 | cmt_trace_exc_o[1];
  assign N224 = N223 | cmt_trace_exc_o[2];
  assign N223 = N222 | cmt_trace_exc_o[3];
  assign N222 = N221 | cmt_trace_exc_o[4];
  assign N221 = cmt_trace_exc_o[6] | cmt_trace_exc_o[5];
  assign calc_status_o[114] = N236 & cmt_trace_stage_reg_o[32];
  assign N236 = cmt_trace_stage_reg_o[34] & N235;
  assign N235 = ~N234;
  assign N234 = N233 | cmt_trace_exc_o[0];
  assign N233 = N232 | cmt_trace_exc_o[1];
  assign N232 = N231 | cmt_trace_exc_o[2];
  assign N231 = N230 | cmt_trace_exc_o[3];
  assign N230 = N229 | cmt_trace_exc_o[4];
  assign N229 = cmt_trace_exc_o[6] | cmt_trace_exc_o[5];
  assign calc_status_o[68] = calc_stage_r_2__decode__pipe_mem_v_ & N243;
  assign N243 = ~N242;
  assign N242 = N241 | exc_stage_r_2__cache_miss_v_;
  assign N241 = N240 | exc_stage_r_2__store_fault_v_;
  assign N240 = N239 | exc_stage_r_2__load_fault_v_;
  assign N239 = N238 | exc_stage_r_2__tlb_miss_v_;
  assign N238 = N237 | exc_stage_r_2__illegal_instr_v_;
  assign N237 = exc_stage_r_2__poison_v_ | exc_stage_r_2__roll_v_;
  assign calc_status_o[3] = N245 & N252;
  assign N245 = exc_stage_n_3__cache_miss_v_ & N244;
  assign N244 = calc_stage_r_2__decode__dcache_r_v_ | calc_stage_r_2__decode__dcache_w_v_;
  assign N252 = ~N251;
  assign N251 = N250 | exc_stage_r_2__cache_miss_v_;
  assign N250 = N249 | exc_stage_r_2__store_fault_v_;
  assign N249 = N248 | exc_stage_r_2__load_fault_v_;
  assign N248 = N247 | exc_stage_r_2__tlb_miss_v_;
  assign N247 = N246 | exc_stage_r_2__illegal_instr_v_;
  assign N246 = exc_stage_r_2__poison_v_ | exc_stage_r_2__roll_v_;
  assign calc_status_o[0] = calc_stage_r_2__decode__instr_v_ & N253;
  assign N253 = ~exc_stage_n_3__roll_v_;
  assign comp_stage_n_slice_iwb_v[1] = calc_stage_r_0__decode__irf_w_v_ & N260;
  assign N260 = ~N259;
  assign N259 = N258 | exc_stage_r_0__cache_miss_v_;
  assign N258 = N257 | exc_stage_r_0__store_fault_v_;
  assign N257 = N256 | exc_stage_r_0__load_fault_v_;
  assign N256 = N255 | exc_stage_r_0__tlb_miss_v_;
  assign N255 = N254 | exc_stage_r_0__illegal_instr_v_;
  assign N254 = exc_stage_r_0__poison_v_ | exc_stage_r_0__roll_v_;
  assign comp_stage_n_slice_fwb_v[1] = calc_stage_r_0__decode__frf_w_v_ & N267;
  assign N267 = ~N266;
  assign N266 = N265 | exc_stage_r_0__cache_miss_v_;
  assign N265 = N264 | exc_stage_r_0__store_fault_v_;
  assign N264 = N263 | exc_stage_r_0__load_fault_v_;
  assign N263 = N262 | exc_stage_r_0__tlb_miss_v_;
  assign N262 = N261 | exc_stage_r_0__illegal_instr_v_;
  assign N261 = exc_stage_r_0__poison_v_ | exc_stage_r_0__roll_v_;
  assign comp_stage_n_slice_iwb_v[2] = calc_stage_r_1__decode__irf_w_v_ & N274;
  assign N274 = ~N273;
  assign N273 = N272 | exc_stage_r_1__cache_miss_v_;
  assign N272 = N271 | exc_stage_r_1__store_fault_v_;
  assign N271 = N270 | exc_stage_r_1__load_fault_v_;
  assign N270 = N269 | exc_stage_r_1__tlb_miss_v_;
  assign N269 = N268 | exc_stage_r_1__illegal_instr_v_;
  assign N268 = exc_stage_r_1__poison_v_ | exc_stage_r_1__roll_v_;
  assign comp_stage_n_slice_fwb_v[2] = calc_stage_r_1__decode__frf_w_v_ & N281;
  assign N281 = ~N280;
  assign N280 = N279 | exc_stage_r_1__cache_miss_v_;
  assign N279 = N278 | exc_stage_r_1__store_fault_v_;
  assign N278 = N277 | exc_stage_r_1__load_fault_v_;
  assign N277 = N276 | exc_stage_r_1__tlb_miss_v_;
  assign N276 = N275 | exc_stage_r_1__illegal_instr_v_;
  assign N275 = exc_stage_r_1__poison_v_ | exc_stage_r_1__roll_v_;
  assign comp_stage_n_slice_iwb_v[3] = calc_stage_r_2__decode__irf_w_v_ & N288;
  assign N288 = ~N287;
  assign N287 = N286 | exc_stage_r_2__cache_miss_v_;
  assign N286 = N285 | exc_stage_r_2__store_fault_v_;
  assign N285 = N284 | exc_stage_r_2__load_fault_v_;
  assign N284 = N283 | exc_stage_r_2__tlb_miss_v_;
  assign N283 = N282 | exc_stage_r_2__illegal_instr_v_;
  assign N282 = exc_stage_r_2__poison_v_ | exc_stage_r_2__roll_v_;
  assign comp_stage_n_slice_fwb_v[3] = calc_stage_r_2__decode__frf_w_v_ & N295;
  assign N295 = ~N294;
  assign N294 = N293 | exc_stage_r_2__cache_miss_v_;
  assign N293 = N292 | exc_stage_r_2__store_fault_v_;
  assign N292 = N291 | exc_stage_r_2__load_fault_v_;
  assign N291 = N290 | exc_stage_r_2__tlb_miss_v_;
  assign N290 = N289 | exc_stage_r_2__illegal_instr_v_;
  assign N289 = exc_stage_r_2__poison_v_ | exc_stage_r_2__roll_v_;
  assign comp_stage_n_slice_iwb_v[4] = calc_stage_r_3__decode__irf_w_v_ & N302;
  assign N302 = ~N301;
  assign N301 = N300 | exc_stage_r_3__cache_miss_v_;
  assign N300 = N299 | exc_stage_r_3__store_fault_v_;
  assign N299 = N298 | exc_stage_r_3__load_fault_v_;
  assign N298 = N297 | exc_stage_r_3__tlb_miss_v_;
  assign N297 = N296 | exc_stage_r_3__illegal_instr_v_;
  assign N296 = exc_stage_r_3__poison_v_ | exc_stage_r_3__roll_v_;
  assign comp_stage_n_slice_fwb_v[4] = calc_stage_r_3__decode__frf_w_v_ & N309;
  assign N309 = ~N308;
  assign N308 = N307 | exc_stage_r_3__cache_miss_v_;
  assign N307 = N306 | exc_stage_r_3__store_fault_v_;
  assign N306 = N305 | exc_stage_r_3__load_fault_v_;
  assign N305 = N304 | exc_stage_r_3__tlb_miss_v_;
  assign N304 = N303 | exc_stage_r_3__illegal_instr_v_;
  assign N303 = exc_stage_r_3__poison_v_ | exc_stage_r_3__roll_v_;
  assign exc_stage_n_1__poison_v_ = exc_stage_r_0__poison_v_ | chk_poison_ex_i;
  assign exc_stage_n_1__roll_v_ = exc_stage_r_0__roll_v_ | chk_roll_i;
  assign exc_stage_n_2__poison_v_ = exc_stage_r_1__poison_v_ | chk_poison_ex_i;
  assign exc_stage_n_2__roll_v_ = exc_stage_r_1__roll_v_ | chk_roll_i;
  assign exc_stage_n_3__roll_v_ = exc_stage_r_2__roll_v_ | chk_roll_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p96_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [95:0] data_i;
  input [5:0] addr_i;
  input [95:0] w_mask_i;
  output [95:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [95:0] data_o;

  hard_mem_1rw_bit_mask_d64_w96_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [8:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  hard_mem_1rw_byte_mask_d512_w64_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_scan_width_p8_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[0] | 1'b0;
  assign t_1__6_ = i[1] | i[0];
  assign t_1__5_ = i[2] | i[1];
  assign t_1__4_ = i[3] | i[2];
  assign t_1__3_ = i[4] | i[3];
  assign t_1__2_ = i[5] | i[4];
  assign t_1__1_ = i[6] | i[5];
  assign t_1__0_ = i[7] | i[6];
  assign t_2__7_ = t_1__7_ | 1'b0;
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__7_ | 1'b0;
  assign o[1] = t_2__6_ | 1'b0;
  assign o[2] = t_2__5_ | 1'b0;
  assign o[3] = t_2__4_ | 1'b0;
  assign o[4] = t_2__3_ | t_2__7_;
  assign o[5] = t_2__2_ | t_2__6_;
  assign o[6] = t_2__1_ | t_2__5_;
  assign o[7] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_width_p8_lo_to_hi_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire N0,N1,N2,N3,N4,N5,N6;
  wire [7:1] scan_lo;

  bsg_scan_width_p8_or_p1_lo_to_hi_p1
  scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[7] = scan_lo[7] & N0;
  assign N0 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N1;
  assign N1 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N2;
  assign N2 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N3;
  assign N3 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N4;
  assign N4 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N5;
  assign N5 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N6;
  assign N6 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_priority_encode_width_p8_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [7:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p8_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_width_p8_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bp_be_dcache_wbuf_queue_width_p97
(
  clk_i,
  data_i,
  el0_en_i,
  el1_en_i,
  mux0_sel_i,
  mux1_sel_i,
  el0_snoop_o,
  el1_snoop_o,
  data_o
);

  input [96:0] data_i;
  output [96:0] el0_snoop_o;
  output [96:0] el1_snoop_o;
  output [96:0] data_o;
  input clk_i;
  input el0_en_i;
  input el1_en_i;
  input mux0_sel_i;
  input mux1_sel_i;
  wire [96:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102;
  reg [96:0] el0_snoop_o,el1_snoop_o;
  assign { N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5 } = (N0)? el0_snoop_o : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N1)? data_i : 1'b0;
  assign N0 = mux0_sel_i;
  assign N1 = N4;
  assign data_o = (N2)? el1_snoop_o : 
                  (N3)? data_i : 1'b0;
  assign N2 = mux1_sel_i;
  assign N3 = N102;
  assign N4 = ~mux0_sel_i;
  assign N102 = ~mux1_sel_i;

  always @(posedge clk_i) begin
    if(el0_en_i) begin
      { el0_snoop_o[96:0] } <= { data_i[96:0] };
    end 
    if(el1_en_i) begin
      { el1_snoop_o[96:0] } <= { N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5 };
    end 
  end


endmodule



module bsg_mux_segmented_segments_p8_segment_width_p8
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [63:0] data0_i;
  input [63:0] data1_i;
  input [7:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;
  assign data_o[7:0] = (N0)? data1_i[7:0] : 
                       (N8)? data0_i[7:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[15:8] = (N1)? data1_i[15:8] : 
                        (N9)? data0_i[15:8] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[23:16] = (N2)? data1_i[23:16] : 
                         (N10)? data0_i[23:16] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[31:24] = (N3)? data1_i[31:24] : 
                         (N11)? data0_i[31:24] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[39:32] = (N4)? data1_i[39:32] : 
                         (N12)? data0_i[39:32] : 1'b0;
  assign N4 = sel_i[4];
  assign data_o[47:40] = (N5)? data1_i[47:40] : 
                         (N13)? data0_i[47:40] : 1'b0;
  assign N5 = sel_i[5];
  assign data_o[55:48] = (N6)? data1_i[55:48] : 
                         (N14)? data0_i[55:48] : 1'b0;
  assign N6 = sel_i[6];
  assign data_o[63:56] = (N7)? data1_i[63:56] : 
                         (N15)? data0_i[63:56] : 1'b0;
  assign N7 = sel_i[7];
  assign N8 = ~sel_i[0];
  assign N9 = ~sel_i[1];
  assign N10 = ~sel_i[2];
  assign N11 = ~sel_i[3];
  assign N12 = ~sel_i[4];
  assign N13 = ~sel_i[5];
  assign N14 = ~sel_i[6];
  assign N15 = ~sel_i[7];

endmodule



module bp_be_dcache_wbuf_data_width_p64_paddr_width_p22_ways_p8_sets_p64
(
  clk_i,
  reset_i,
  v_i,
  wbuf_entry_i,
  yumi_i,
  v_o,
  wbuf_entry_o,
  empty_o,
  bypass_addr_i,
  bypass_v_i,
  bypass_data_o,
  bypass_mask_o,
  lce_snoop_index_i,
  lce_snoop_way_i,
  lce_snoop_match_o
);

  input [96:0] wbuf_entry_i;
  output [96:0] wbuf_entry_o;
  input [21:0] bypass_addr_i;
  output [63:0] bypass_data_o;
  output [7:0] bypass_mask_o;
  input [5:0] lce_snoop_index_i;
  input [2:0] lce_snoop_way_i;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input bypass_v_i;
  output v_o;
  output empty_o;
  output lce_snoop_match_o;
  wire [96:0] wbuf_entry_o,wbuf_entry_el0,wbuf_entry_el1;
  wire v_o,empty_o,lce_snoop_match_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  el0_valid,el1_valid,el0_enable,N14,el1_enable,mux0_sel,mux1_sel,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,tag_hit0_n,tag_hit1_n,tag_hit2_n,n_2_net__7_,
  n_2_net__6_,n_2_net__5_,n_2_net__4_,n_2_net__3_,n_2_net__2_,n_2_net__1_,n_2_net__0_,
  n_4_net__7_,n_4_net__6_,n_4_net__5_,n_4_net__4_,n_4_net__3_,n_4_net__2_,n_4_net__1_,
  n_4_net__0_,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,
  N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,lce_snoop_el2_match,N105,N106,lce_snoop_el0_match,N107,N108,
  lce_snoop_el1_match,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,
  N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
  N139,N140,N141,N142,N143,N144,N145;
  wire [7:7] tag_hit0x4,tag_hit1x4,tag_hit2x4;
  wire [7:0] bypass_mask_n;
  wire [63:0] el0or1_data,bypass_data_n;
  reg [1:0] num_els_r;
  reg [63:0] bypass_data_o;
  reg [7:0] bypass_mask_o;
  assign N8 = N6 & N7;
  assign N9 = num_els_r[1] | N7;
  assign N11 = N6 | num_els_r[0];
  assign N13 = num_els_r[1] & num_els_r[0];

  bp_be_dcache_wbuf_queue_width_p97
  wbq
  (
    .clk_i(clk_i),
    .data_i(wbuf_entry_i),
    .el0_en_i(el0_enable),
    .el1_en_i(el1_enable),
    .mux0_sel_i(mux0_sel),
    .mux1_sel_i(mux1_sel),
    .el0_snoop_o(wbuf_entry_el0),
    .el1_snoop_o(wbuf_entry_el1),
    .data_o(wbuf_entry_o)
  );

  assign tag_hit0_n = bypass_addr_i[21:3] == wbuf_entry_el0[96:78];
  assign tag_hit1_n = bypass_addr_i[21:3] == wbuf_entry_el1[96:78];
  assign tag_hit2_n = bypass_addr_i[21:3] == wbuf_entry_i[96:78];

  bsg_mux_segmented_segments_p8_segment_width_p8
  mux_segmented_merge0
  (
    .data0_i(wbuf_entry_el1[74:11]),
    .data1_i(wbuf_entry_el0[74:11]),
    .sel_i({ n_2_net__7_, n_2_net__6_, n_2_net__5_, n_2_net__4_, n_2_net__3_, n_2_net__2_, n_2_net__1_, n_2_net__0_ }),
    .data_o(el0or1_data)
  );


  bsg_mux_segmented_segments_p8_segment_width_p8
  mux_segmented_merge1
  (
    .data0_i(el0or1_data),
    .data1_i(wbuf_entry_i[74:11]),
    .sel_i({ n_4_net__7_, n_4_net__6_, n_4_net__5_, n_4_net__4_, n_4_net__3_, n_4_net__2_, n_4_net__1_, n_4_net__0_ }),
    .data_o(bypass_data_n)
  );

  assign N103 = lce_snoop_index_i == wbuf_entry_i[86:81];
  assign N104 = lce_snoop_way_i == wbuf_entry_i[2:0];
  assign N105 = lce_snoop_index_i == wbuf_entry_el0[86:81];
  assign N106 = lce_snoop_way_i == wbuf_entry_el0[2:0];
  assign N107 = lce_snoop_index_i == wbuf_entry_el1[86:81];
  assign N108 = lce_snoop_way_i == wbuf_entry_el1[2:0];
  assign { N21, N20 } = v_i - N19;
  assign { N23, N22 } = num_els_r + { N21, N20 };
  assign v_o = (N0)? v_i : 
               (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N8;
  assign N1 = N10;
  assign N2 = N12;
  assign N3 = N13;
  assign empty_o = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b0 : 1'b0;
  assign el0_valid = (N0)? 1'b0 : 
                     (N1)? 1'b0 : 
                     (N2)? 1'b1 : 
                     (N3)? 1'b0 : 1'b0;
  assign el1_valid = (N0)? 1'b0 : 
                     (N1)? 1'b1 : 
                     (N2)? 1'b1 : 
                     (N3)? 1'b0 : 1'b0;
  assign el0_enable = (N0)? 1'b0 : 
                      (N1)? N15 : 
                      (N2)? N17 : 
                      (N3)? 1'b0 : 1'b0;
  assign el1_enable = (N0)? N14 : 
                      (N1)? N16 : 
                      (N2)? yumi_i : 
                      (N3)? 1'b0 : 1'b0;
  assign mux0_sel = (N0)? 1'b0 : 
                    (N1)? 1'b0 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign mux1_sel = (N0)? 1'b0 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign { N25, N24 } = (N4)? { 1'b0, 1'b0 } : 
                        (N5)? { N23, N22 } : 1'b0;
  assign N4 = reset_i;
  assign N5 = N18;
  assign N28 = (N4)? 1'b1 : 
               (N102)? 1'b1 : 
               (N27)? 1'b0 : 1'b0;
  assign { N36, N35, N34, N33, N32, N31, N30, N29 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N102)? bypass_mask_n : 1'b0;
  assign { N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                               (N102)? bypass_data_n : 1'b0;
  assign N6 = ~num_els_r[1];
  assign N7 = ~num_els_r[0];
  assign N10 = ~N9;
  assign N12 = ~N11;
  assign N14 = v_i & N109;
  assign N109 = ~yumi_i;
  assign N15 = v_i & N109;
  assign N16 = v_i & yumi_i;
  assign N17 = v_i & yumi_i;
  assign N18 = ~reset_i;
  assign N19 = v_o & yumi_i;
  assign tag_hit0x4[7] = tag_hit0_n & el0_valid;
  assign tag_hit1x4[7] = tag_hit1_n & el1_valid;
  assign tag_hit2x4[7] = tag_hit2_n & v_i;
  assign bypass_mask_n[7] = N112 | N113;
  assign N112 = N110 | N111;
  assign N110 = tag_hit0x4[7] & wbuf_entry_el0[10];
  assign N111 = tag_hit1x4[7] & wbuf_entry_el1[10];
  assign N113 = tag_hit2x4[7] & wbuf_entry_i[10];
  assign bypass_mask_n[6] = N116 | N117;
  assign N116 = N114 | N115;
  assign N114 = tag_hit0x4[7] & wbuf_entry_el0[9];
  assign N115 = tag_hit1x4[7] & wbuf_entry_el1[9];
  assign N117 = tag_hit2x4[7] & wbuf_entry_i[9];
  assign bypass_mask_n[5] = N120 | N121;
  assign N120 = N118 | N119;
  assign N118 = tag_hit0x4[7] & wbuf_entry_el0[8];
  assign N119 = tag_hit1x4[7] & wbuf_entry_el1[8];
  assign N121 = tag_hit2x4[7] & wbuf_entry_i[8];
  assign bypass_mask_n[4] = N124 | N125;
  assign N124 = N122 | N123;
  assign N122 = tag_hit0x4[7] & wbuf_entry_el0[7];
  assign N123 = tag_hit1x4[7] & wbuf_entry_el1[7];
  assign N125 = tag_hit2x4[7] & wbuf_entry_i[7];
  assign bypass_mask_n[3] = N128 | N129;
  assign N128 = N126 | N127;
  assign N126 = tag_hit0x4[7] & wbuf_entry_el0[6];
  assign N127 = tag_hit1x4[7] & wbuf_entry_el1[6];
  assign N129 = tag_hit2x4[7] & wbuf_entry_i[6];
  assign bypass_mask_n[2] = N132 | N133;
  assign N132 = N130 | N131;
  assign N130 = tag_hit0x4[7] & wbuf_entry_el0[5];
  assign N131 = tag_hit1x4[7] & wbuf_entry_el1[5];
  assign N133 = tag_hit2x4[7] & wbuf_entry_i[5];
  assign bypass_mask_n[1] = N136 | N137;
  assign N136 = N134 | N135;
  assign N134 = tag_hit0x4[7] & wbuf_entry_el0[4];
  assign N135 = tag_hit1x4[7] & wbuf_entry_el1[4];
  assign N137 = tag_hit2x4[7] & wbuf_entry_i[4];
  assign bypass_mask_n[0] = N140 | N141;
  assign N140 = N138 | N139;
  assign N138 = tag_hit0x4[7] & wbuf_entry_el0[3];
  assign N139 = tag_hit1x4[7] & wbuf_entry_el1[3];
  assign N141 = tag_hit2x4[7] & wbuf_entry_i[3];
  assign n_2_net__7_ = tag_hit0x4[7] & wbuf_entry_el0[10];
  assign n_2_net__6_ = tag_hit0x4[7] & wbuf_entry_el0[9];
  assign n_2_net__5_ = tag_hit0x4[7] & wbuf_entry_el0[8];
  assign n_2_net__4_ = tag_hit0x4[7] & wbuf_entry_el0[7];
  assign n_2_net__3_ = tag_hit0x4[7] & wbuf_entry_el0[6];
  assign n_2_net__2_ = tag_hit0x4[7] & wbuf_entry_el0[5];
  assign n_2_net__1_ = tag_hit0x4[7] & wbuf_entry_el0[4];
  assign n_2_net__0_ = tag_hit0x4[7] & wbuf_entry_el0[3];
  assign n_4_net__7_ = tag_hit2x4[7] & wbuf_entry_i[10];
  assign n_4_net__6_ = tag_hit2x4[7] & wbuf_entry_i[9];
  assign n_4_net__5_ = tag_hit2x4[7] & wbuf_entry_i[8];
  assign n_4_net__4_ = tag_hit2x4[7] & wbuf_entry_i[7];
  assign n_4_net__3_ = tag_hit2x4[7] & wbuf_entry_i[6];
  assign n_4_net__2_ = tag_hit2x4[7] & wbuf_entry_i[5];
  assign n_4_net__1_ = tag_hit2x4[7] & wbuf_entry_i[4];
  assign n_4_net__0_ = tag_hit2x4[7] & wbuf_entry_i[3];
  assign N26 = bypass_v_i | reset_i;
  assign N27 = ~N26;
  assign N101 = ~reset_i;
  assign N102 = bypass_v_i & N101;
  assign lce_snoop_el2_match = N142 & N104;
  assign N142 = v_i & N103;
  assign lce_snoop_el0_match = N143 & N106;
  assign N143 = el0_valid & N105;
  assign lce_snoop_el1_match = N144 & N108;
  assign N144 = el1_valid & N107;
  assign lce_snoop_match_o = N145 | lce_snoop_el1_match;
  assign N145 = lce_snoop_el2_match | lce_snoop_el0_match;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { num_els_r[1:0] } <= { N25, N24 };
    end 
    if(N28) begin
      { bypass_data_o[63:0] } <= { N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37 };
      { bypass_mask_o[7:0] } <= { N36, N35, N34, N33, N32, N31, N30, N29 };
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p15_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [14:0] data_i;
  input [5:0] addr_i;
  input [14:0] w_mask_i;
  output [14:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [14:0] data_o;

  hard_mem_1rw_bit_mask_d64_w15_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bp_be_dcache_lru_encode_ways_p8
(
  lru_i,
  way_id_o
);

  input [6:0] lru_i;
  output [2:0] way_id_o;
  wire [2:0] way_id_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30;
  assign N11 = N8 & N9;
  assign N12 = N11 & N10;
  assign N13 = lru_i[3] & N9;
  assign N14 = N13 & N10;
  assign N16 = N15 & lru_i[1];
  assign N17 = N16 & N10;
  assign N18 = lru_i[4] & lru_i[1];
  assign N19 = N18 & N10;
  assign N22 = N20 & N21;
  assign N23 = N22 & lru_i[0];
  assign N24 = lru_i[5] & N21;
  assign N25 = N24 & lru_i[0];
  assign N27 = N26 & lru_i[2];
  assign N28 = N27 & lru_i[0];
  assign N29 = lru_i[6] & lru_i[2];
  assign N30 = N29 & lru_i[0];
  assign way_id_o = (N0)? { 1'b0, 1'b0, 1'b0 } : 
                    (N1)? { 1'b0, 1'b0, 1'b1 } : 
                    (N2)? { 1'b0, 1'b1, 1'b0 } : 
                    (N3)? { 1'b0, 1'b1, 1'b1 } : 
                    (N4)? { 1'b1, 1'b0, 1'b0 } : 
                    (N5)? { 1'b1, 1'b0, 1'b1 } : 
                    (N6)? { 1'b1, 1'b1, 1'b0 } : 
                    (N7)? { 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N0 = N12;
  assign N1 = N14;
  assign N2 = N17;
  assign N3 = N19;
  assign N4 = N23;
  assign N5 = N25;
  assign N6 = N28;
  assign N7 = N30;
  assign N8 = ~lru_i[3];
  assign N9 = ~lru_i[1];
  assign N10 = ~lru_i[0];
  assign N15 = ~lru_i[4];
  assign N20 = ~lru_i[5];
  assign N21 = ~lru_i[2];
  assign N26 = ~lru_i[6];

endmodule



module bp_be_dcache_lce_req_data_width_p64_paddr_width_p22_num_cce_p1_num_lce_p2_ways_p8_sets_p64
(
  clk_i,
  reset_i,
  lce_id_i,
  load_miss_i,
  store_miss_i,
  miss_addr_i,
  lru_way_i,
  dirty_i,
  cache_miss_o,
  tr_received_i,
  cce_data_received_i,
  tag_set_i,
  tag_set_wakeup_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i
);

  input [0:0] lce_id_i;
  input [21:0] miss_addr_i;
  input [2:0] lru_way_i;
  input [7:0] dirty_i;
  output [29:0] lce_req_o;
  output [25:0] lce_resp_o;
  input clk_i;
  input reset_i;
  input load_miss_i;
  input store_miss_i;
  input tr_received_i;
  input cce_data_received_i;
  input tag_set_i;
  input tag_set_wakeup_i;
  input lce_req_ready_i;
  input lce_resp_yumi_i;
  output cache_miss_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  wire [25:0] lce_resp_o;
  wire cache_miss_o,lce_req_v_o,lce_resp_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,missed,
  tr_received,cce_data_received,tag_set,dirty_lru_flopped_n,tr_received_n,
  cce_data_received_n,tag_set_n,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,
  N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,
  N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,
  N120,N121,N122,N123,N124;
  wire [2:0] state_n;
  reg [29:0] lce_req_o;
  reg [2:0] state_r,lru_way_r;
  reg dirty_lru_flopped_r,tr_received_r,cce_data_received_r,tag_set_r,
  load_not_store_r,dirty_r;
  assign lce_resp_o[23] = 1'b1;
  assign lce_resp_o[25] = 1'b0;
  assign lce_req_o[26] = 1'b0;
  assign lce_req_o[29] = 1'b0;
  assign lce_resp_o[21] = lce_req_o[25];
  assign lce_resp_o[20] = lce_req_o[24];
  assign lce_resp_o[19] = lce_req_o[23];
  assign lce_resp_o[18] = lce_req_o[22];
  assign lce_resp_o[17] = lce_req_o[21];
  assign lce_resp_o[16] = lce_req_o[20];
  assign lce_resp_o[15] = lce_req_o[19];
  assign lce_resp_o[14] = lce_req_o[18];
  assign lce_resp_o[13] = lce_req_o[17];
  assign lce_resp_o[12] = lce_req_o[16];
  assign lce_resp_o[11] = lce_req_o[15];
  assign lce_resp_o[10] = lce_req_o[14];
  assign lce_resp_o[9] = lce_req_o[13];
  assign lce_resp_o[8] = lce_req_o[12];
  assign lce_resp_o[7] = lce_req_o[11];
  assign lce_resp_o[6] = lce_req_o[10];
  assign lce_resp_o[5] = lce_req_o[9];
  assign lce_resp_o[4] = lce_req_o[8];
  assign lce_resp_o[3] = lce_req_o[7];
  assign lce_resp_o[2] = lce_req_o[6];
  assign lce_resp_o[1] = lce_req_o[5];
  assign lce_resp_o[0] = lce_req_o[4];
  assign lce_resp_o[24] = lce_id_i[0];
  assign lce_req_o[28] = lce_id_i[0];
  assign N27 = (N19)? dirty_i[0] : 
               (N21)? dirty_i[1] : 
               (N23)? dirty_i[2] : 
               (N25)? dirty_i[3] : 
               (N20)? dirty_i[4] : 
               (N22)? dirty_i[5] : 
               (N24)? dirty_i[6] : 
               (N26)? dirty_i[7] : 1'b0;
  assign N31 = N28 & N29;
  assign N32 = N31 & N30;
  assign N33 = state_r[2] | state_r[1];
  assign N34 = N33 | N30;
  assign N36 = N28 | state_r[1];
  assign N37 = N36 | state_r[0];
  assign N39 = state_r[2] | N29;
  assign N40 = N39 | state_r[0];
  assign N42 = state_r[2] | N29;
  assign N43 = N42 | N30;
  assign N45 = state_r[2] & state_r[0];
  assign N46 = state_r[2] & state_r[1];
  assign lce_req_o[3:1] = (N0)? lru_way_r : 
                          (N1)? lru_way_i : 1'b0;
  assign N0 = dirty_lru_flopped_r;
  assign N1 = N11;
  assign lce_req_o[0] = (N0)? dirty_r : 
                        (N1)? N27 : 1'b0;
  assign { N59, N58, N57 } = (N2)? { 1'b0, 1'b1, 1'b0 } : 
                             (N67)? { 1'b0, 1'b1, 1'b1 } : 
                             (N56)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N2 = tr_received;
  assign { N62, N61, N60 } = (N3)? { 1'b0, 1'b0, 1'b0 } : 
                             (N65)? { N59, N58, N57 } : 
                             (N54)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N3 = tag_set_wakeup_i;
  assign cache_miss_o = (N4)? missed : 
                        (N5)? 1'b1 : 
                        (N6)? 1'b1 : 
                        (N7)? 1'b1 : 
                        (N8)? 1'b1 : 
                        (N9)? 1'b0 : 1'b0;
  assign N4 = N32;
  assign N5 = N35;
  assign N6 = N38;
  assign N7 = N41;
  assign N8 = N44;
  assign N9 = N47;
  assign state_n = (N4)? { 1'b0, 1'b0, 1'b1 } : 
                   (N5)? { lce_req_ready_i, 1'b0, N49 } : 
                   (N6)? { N62, N61, N60 } : 
                   (N7)? { 1'b0, N63, 1'b0 } : 
                   (N8)? { 1'b0, N63, N63 } : 
                   (N9)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign dirty_lru_flopped_n = (N4)? 1'b0 : 
                               (N5)? 1'b1 : 1'b0;
  assign tr_received_n = (N4)? 1'b0 : 
                         (N6)? 1'b1 : 1'b0;
  assign cce_data_received_n = (N4)? 1'b0 : 
                               (N6)? 1'b1 : 1'b0;
  assign tag_set_n = (N4)? 1'b0 : 
                     (N6)? 1'b1 : 1'b0;
  assign lce_req_v_o = (N4)? 1'b0 : 
                       (N5)? 1'b1 : 
                       (N6)? 1'b0 : 
                       (N7)? 1'b0 : 
                       (N8)? 1'b0 : 
                       (N9)? 1'b0 : 1'b0;
  assign lce_resp_v_o = (N4)? 1'b0 : 
                        (N5)? 1'b0 : 
                        (N6)? 1'b0 : 
                        (N7)? 1'b1 : 
                        (N8)? 1'b1 : 
                        (N9)? 1'b0 : 1'b0;
  assign lce_resp_o[22] = (N4)? 1'b0 : 
                          (N5)? 1'b0 : 
                          (N6)? 1'b0 : 
                          (N7)? 1'b0 : 
                          (N8)? 1'b1 : 
                          (N9)? 1'b0 : 1'b0;
  assign missed = load_miss_i | store_miss_i;
  assign tr_received = tr_received_r | tr_received_i;
  assign cce_data_received = cce_data_received_r | cce_data_received_i;
  assign tag_set = tag_set_r | tag_set_i;
  assign N10 = ~load_not_store_r;
  assign lce_req_o[27] = N10;
  assign N11 = ~dirty_lru_flopped_r;
  assign N12 = ~lru_way_i[0];
  assign N13 = ~lru_way_i[1];
  assign N14 = N12 & N13;
  assign N15 = N12 & lru_way_i[1];
  assign N16 = lru_way_i[0] & N13;
  assign N17 = lru_way_i[0] & lru_way_i[1];
  assign N18 = ~lru_way_i[2];
  assign N19 = N14 & N18;
  assign N20 = N14 & lru_way_i[2];
  assign N21 = N16 & N18;
  assign N22 = N16 & lru_way_i[2];
  assign N23 = N15 & N18;
  assign N24 = N15 & lru_way_i[2];
  assign N25 = N17 & N18;
  assign N26 = N17 & lru_way_i[2];
  assign N28 = ~state_r[2];
  assign N29 = ~state_r[1];
  assign N30 = ~state_r[0];
  assign N35 = ~N34;
  assign N38 = ~N37;
  assign N41 = ~N40;
  assign N44 = ~N43;
  assign N47 = N45 | N46;
  assign N48 = ~missed;
  assign N49 = ~lce_req_ready_i;
  assign N50 = ~tr_received_i;
  assign N51 = ~cce_data_received_i;
  assign N52 = ~tag_set_i;
  assign N53 = tag_set | tag_set_wakeup_i;
  assign N54 = ~N53;
  assign N55 = cce_data_received | tr_received;
  assign N56 = ~N55;
  assign N63 = ~lce_resp_yumi_i;
  assign N64 = ~tag_set_wakeup_i;
  assign N65 = tag_set & N64;
  assign N66 = ~tr_received;
  assign N67 = cce_data_received & N66;
  assign N68 = ~reset_i;
  assign N69 = N32 & N68;
  assign N70 = N48 & N69;
  assign N71 = N35 & N68;
  assign N72 = N70 | N71;
  assign N73 = N38 & N68;
  assign N74 = N72 | N73;
  assign N75 = N41 & N68;
  assign N76 = N74 | N75;
  assign N77 = N44 & N68;
  assign N78 = N76 | N77;
  assign N79 = N47 & N68;
  assign N80 = N78 | N79;
  assign N81 = ~N80;
  assign N82 = N68 & N81;
  assign N83 = N48 & N32;
  assign N84 = ~N83;
  assign N85 = N83 | N38;
  assign N86 = N85 | N41;
  assign N87 = N86 | N44;
  assign N88 = N87 | N47;
  assign N89 = ~N88;
  assign N90 = N83 | N35;
  assign N91 = N50 & N38;
  assign N92 = N90 | N91;
  assign N93 = N92 | N41;
  assign N94 = N93 | N44;
  assign N95 = N94 | N47;
  assign N96 = ~N95;
  assign N97 = N51 & N38;
  assign N98 = N90 | N97;
  assign N99 = N98 | N41;
  assign N100 = N99 | N44;
  assign N101 = N100 | N47;
  assign N102 = ~N101;
  assign N103 = N52 & N38;
  assign N104 = N90 | N103;
  assign N105 = N104 | N41;
  assign N106 = N105 | N44;
  assign N107 = N106 | N47;
  assign N108 = ~N107;
  assign N109 = dirty_lru_flopped_r & N71;
  assign N110 = N69 | N109;
  assign N111 = N110 | N73;
  assign N112 = N111 | N75;
  assign N113 = N112 | N77;
  assign N114 = N113 | N79;
  assign N115 = ~N114;
  assign N116 = N68 & N115;
  assign N117 = dirty_lru_flopped_r & N71;
  assign N118 = N69 | N117;
  assign N119 = N118 | N73;
  assign N120 = N119 | N75;
  assign N121 = N120 | N77;
  assign N122 = N121 | N79;
  assign N123 = ~N122;
  assign N124 = N68 & N123;

  always @(posedge clk_i) begin
    if(N82) begin
      { lce_req_o[25:4] } <= { miss_addr_i[21:0] };
      load_not_store_r <= load_miss_i;
    end 
    if(reset_i) begin
      { state_r[2:0] } <= { 1'b0, 1'b0, 1'b0 };
    end else if(N84) begin
      { state_r[2:0] } <= { state_n[2:0] };
    end 
    if(reset_i) begin
      dirty_lru_flopped_r <= 1'b0;
    end else if(N89) begin
      dirty_lru_flopped_r <= dirty_lru_flopped_n;
    end 
    if(reset_i) begin
      tr_received_r <= 1'b0;
    end else if(N96) begin
      tr_received_r <= tr_received_n;
    end 
    if(reset_i) begin
      cce_data_received_r <= 1'b0;
    end else if(N102) begin
      cce_data_received_r <= cce_data_received_n;
    end 
    if(reset_i) begin
      tag_set_r <= 1'b0;
    end else if(N108) begin
      tag_set_r <= tag_set_n;
    end 
    if(N116) begin
      { lru_way_r[2:0] } <= { lru_way_i[2:0] };
    end 
    if(N124) begin
      dirty_r <= N27;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p36_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [35:0] w_data_i;
  input [0:0] r_addr_i;
  output [35:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [35:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [71:0] mem;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[71] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[70] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[69] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[68] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[67] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[66] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[65] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[64] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[63] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[62] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[61] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[60] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[59] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[58] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[57] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[56] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[55] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[54] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[53] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[52] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[51] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[47] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[46] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[45] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[44] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[43] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[42] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[41] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[40] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[39] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[38] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[37] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[36] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[71:36] } <= { w_data_i[35:0] };
    end 
    if(N7) begin
      { mem[35:0] } <= { w_data_i[35:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p36_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [35:0] w_data_i;
  input [0:0] r_addr_i;
  output [35:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [35:0] r_data_o;

  bsg_mem_1r1w_synth_width_p36_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p36
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [35:0] data_i;
  output [35:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [35:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p36_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bp_be_dcache_lce_cmd_num_cce_p1_num_lce_p2_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_data_width_p64
(
  clk_i,
  reset_i,
  lce_id_i,
  lce_sync_done_o,
  tag_set_o,
  tag_set_wakeup_o,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_yumi_o,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_tr_resp_o,
  lce_tr_resp_v_o,
  lce_tr_resp_ready_i,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_data_i,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_v_o,
  tag_mem_pkt_o,
  tag_mem_pkt_yumi_i,
  stat_mem_pkt_v_o,
  stat_mem_pkt_o,
  dirty_i,
  stat_mem_pkt_yumi_i
);

  input [0:0] lce_id_i;
  input [35:0] lce_cmd_i;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  output [538:0] lce_tr_resp_o;
  output [521:0] data_mem_pkt_o;
  input [511:0] data_mem_data_i;
  output [22:0] tag_mem_pkt_o;
  output [10:0] stat_mem_pkt_o;
  input [7:0] dirty_i;
  input clk_i;
  input reset_i;
  input lce_cmd_v_i;
  input lce_resp_yumi_i;
  input lce_data_resp_ready_i;
  input lce_tr_resp_ready_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input stat_mem_pkt_yumi_i;
  output lce_sync_done_o;
  output tag_set_o;
  output tag_set_wakeup_o;
  output lce_cmd_yumi_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_tr_resp_v_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output stat_mem_pkt_v_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [538:0] lce_tr_resp_o;
  wire [521:0] data_mem_pkt_o;
  wire [22:0] tag_mem_pkt_o;
  wire [10:0] stat_mem_pkt_o;
  wire lce_sync_done_o,tag_set_o,tag_set_wakeup_o,lce_cmd_yumi_o,lce_resp_v_o,
  lce_data_resp_v_o,lce_tr_resp_v_o,data_mem_pkt_v_o,tag_mem_pkt_v_o,stat_mem_pkt_v_o,N0,
  N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,lce_tr_resp_done,lce_data_resp_done,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,
  N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
  N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,
  N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,
  N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,
  N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
  N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,
  N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,
  N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,
  N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,
  N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,
  N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,
  N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,
  N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,
  N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,
  N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,
  N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,
  N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,
  N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
  N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,
  N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,
  N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,
  N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,
  N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,
  N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
  N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,
  N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,
  N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,
  N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,
  N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,
  N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,
  N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1606,
  N1607;
  wire [2:0] state_n;
  reg [511:0] data_buf_r;
  reg [2:0] state_r;
  reg [0:0] sync_ack_count_r;
  reg tr_data_buffered_r,wb_data_buffered_r,wb_data_read_r,wb_dirty_cleared_r,
  invalidated_tag_r;
  assign data_mem_pkt_o[0] = 1'b0;
  assign data_mem_pkt_o[1] = 1'b0;
  assign data_mem_pkt_o[2] = 1'b0;
  assign data_mem_pkt_o[3] = 1'b0;
  assign data_mem_pkt_o[4] = 1'b0;
  assign data_mem_pkt_o[5] = 1'b0;
  assign data_mem_pkt_o[6] = 1'b0;
  assign data_mem_pkt_o[7] = 1'b0;
  assign data_mem_pkt_o[8] = 1'b0;
  assign data_mem_pkt_o[9] = 1'b0;
  assign data_mem_pkt_o[10] = 1'b0;
  assign data_mem_pkt_o[11] = 1'b0;
  assign data_mem_pkt_o[12] = 1'b0;
  assign data_mem_pkt_o[13] = 1'b0;
  assign data_mem_pkt_o[14] = 1'b0;
  assign data_mem_pkt_o[15] = 1'b0;
  assign data_mem_pkt_o[16] = 1'b0;
  assign data_mem_pkt_o[17] = 1'b0;
  assign data_mem_pkt_o[18] = 1'b0;
  assign data_mem_pkt_o[19] = 1'b0;
  assign data_mem_pkt_o[20] = 1'b0;
  assign data_mem_pkt_o[21] = 1'b0;
  assign data_mem_pkt_o[22] = 1'b0;
  assign data_mem_pkt_o[23] = 1'b0;
  assign data_mem_pkt_o[24] = 1'b0;
  assign data_mem_pkt_o[25] = 1'b0;
  assign data_mem_pkt_o[26] = 1'b0;
  assign data_mem_pkt_o[27] = 1'b0;
  assign data_mem_pkt_o[28] = 1'b0;
  assign data_mem_pkt_o[29] = 1'b0;
  assign data_mem_pkt_o[30] = 1'b0;
  assign data_mem_pkt_o[31] = 1'b0;
  assign data_mem_pkt_o[32] = 1'b0;
  assign data_mem_pkt_o[33] = 1'b0;
  assign data_mem_pkt_o[34] = 1'b0;
  assign data_mem_pkt_o[35] = 1'b0;
  assign data_mem_pkt_o[36] = 1'b0;
  assign data_mem_pkt_o[37] = 1'b0;
  assign data_mem_pkt_o[38] = 1'b0;
  assign data_mem_pkt_o[39] = 1'b0;
  assign data_mem_pkt_o[40] = 1'b0;
  assign data_mem_pkt_o[41] = 1'b0;
  assign data_mem_pkt_o[42] = 1'b0;
  assign data_mem_pkt_o[43] = 1'b0;
  assign data_mem_pkt_o[44] = 1'b0;
  assign data_mem_pkt_o[45] = 1'b0;
  assign data_mem_pkt_o[46] = 1'b0;
  assign data_mem_pkt_o[47] = 1'b0;
  assign data_mem_pkt_o[48] = 1'b0;
  assign data_mem_pkt_o[49] = 1'b0;
  assign data_mem_pkt_o[50] = 1'b0;
  assign data_mem_pkt_o[51] = 1'b0;
  assign data_mem_pkt_o[52] = 1'b0;
  assign data_mem_pkt_o[53] = 1'b0;
  assign data_mem_pkt_o[54] = 1'b0;
  assign data_mem_pkt_o[55] = 1'b0;
  assign data_mem_pkt_o[56] = 1'b0;
  assign data_mem_pkt_o[57] = 1'b0;
  assign data_mem_pkt_o[58] = 1'b0;
  assign data_mem_pkt_o[59] = 1'b0;
  assign data_mem_pkt_o[60] = 1'b0;
  assign data_mem_pkt_o[61] = 1'b0;
  assign data_mem_pkt_o[62] = 1'b0;
  assign data_mem_pkt_o[63] = 1'b0;
  assign data_mem_pkt_o[64] = 1'b0;
  assign data_mem_pkt_o[65] = 1'b0;
  assign data_mem_pkt_o[66] = 1'b0;
  assign data_mem_pkt_o[67] = 1'b0;
  assign data_mem_pkt_o[68] = 1'b0;
  assign data_mem_pkt_o[69] = 1'b0;
  assign data_mem_pkt_o[70] = 1'b0;
  assign data_mem_pkt_o[71] = 1'b0;
  assign data_mem_pkt_o[72] = 1'b0;
  assign data_mem_pkt_o[73] = 1'b0;
  assign data_mem_pkt_o[74] = 1'b0;
  assign data_mem_pkt_o[75] = 1'b0;
  assign data_mem_pkt_o[76] = 1'b0;
  assign data_mem_pkt_o[77] = 1'b0;
  assign data_mem_pkt_o[78] = 1'b0;
  assign data_mem_pkt_o[79] = 1'b0;
  assign data_mem_pkt_o[80] = 1'b0;
  assign data_mem_pkt_o[81] = 1'b0;
  assign data_mem_pkt_o[82] = 1'b0;
  assign data_mem_pkt_o[83] = 1'b0;
  assign data_mem_pkt_o[84] = 1'b0;
  assign data_mem_pkt_o[85] = 1'b0;
  assign data_mem_pkt_o[86] = 1'b0;
  assign data_mem_pkt_o[87] = 1'b0;
  assign data_mem_pkt_o[88] = 1'b0;
  assign data_mem_pkt_o[89] = 1'b0;
  assign data_mem_pkt_o[90] = 1'b0;
  assign data_mem_pkt_o[91] = 1'b0;
  assign data_mem_pkt_o[92] = 1'b0;
  assign data_mem_pkt_o[93] = 1'b0;
  assign data_mem_pkt_o[94] = 1'b0;
  assign data_mem_pkt_o[95] = 1'b0;
  assign data_mem_pkt_o[96] = 1'b0;
  assign data_mem_pkt_o[97] = 1'b0;
  assign data_mem_pkt_o[98] = 1'b0;
  assign data_mem_pkt_o[99] = 1'b0;
  assign data_mem_pkt_o[100] = 1'b0;
  assign data_mem_pkt_o[101] = 1'b0;
  assign data_mem_pkt_o[102] = 1'b0;
  assign data_mem_pkt_o[103] = 1'b0;
  assign data_mem_pkt_o[104] = 1'b0;
  assign data_mem_pkt_o[105] = 1'b0;
  assign data_mem_pkt_o[106] = 1'b0;
  assign data_mem_pkt_o[107] = 1'b0;
  assign data_mem_pkt_o[108] = 1'b0;
  assign data_mem_pkt_o[109] = 1'b0;
  assign data_mem_pkt_o[110] = 1'b0;
  assign data_mem_pkt_o[111] = 1'b0;
  assign data_mem_pkt_o[112] = 1'b0;
  assign data_mem_pkt_o[113] = 1'b0;
  assign data_mem_pkt_o[114] = 1'b0;
  assign data_mem_pkt_o[115] = 1'b0;
  assign data_mem_pkt_o[116] = 1'b0;
  assign data_mem_pkt_o[117] = 1'b0;
  assign data_mem_pkt_o[118] = 1'b0;
  assign data_mem_pkt_o[119] = 1'b0;
  assign data_mem_pkt_o[120] = 1'b0;
  assign data_mem_pkt_o[121] = 1'b0;
  assign data_mem_pkt_o[122] = 1'b0;
  assign data_mem_pkt_o[123] = 1'b0;
  assign data_mem_pkt_o[124] = 1'b0;
  assign data_mem_pkt_o[125] = 1'b0;
  assign data_mem_pkt_o[126] = 1'b0;
  assign data_mem_pkt_o[127] = 1'b0;
  assign data_mem_pkt_o[128] = 1'b0;
  assign data_mem_pkt_o[129] = 1'b0;
  assign data_mem_pkt_o[130] = 1'b0;
  assign data_mem_pkt_o[131] = 1'b0;
  assign data_mem_pkt_o[132] = 1'b0;
  assign data_mem_pkt_o[133] = 1'b0;
  assign data_mem_pkt_o[134] = 1'b0;
  assign data_mem_pkt_o[135] = 1'b0;
  assign data_mem_pkt_o[136] = 1'b0;
  assign data_mem_pkt_o[137] = 1'b0;
  assign data_mem_pkt_o[138] = 1'b0;
  assign data_mem_pkt_o[139] = 1'b0;
  assign data_mem_pkt_o[140] = 1'b0;
  assign data_mem_pkt_o[141] = 1'b0;
  assign data_mem_pkt_o[142] = 1'b0;
  assign data_mem_pkt_o[143] = 1'b0;
  assign data_mem_pkt_o[144] = 1'b0;
  assign data_mem_pkt_o[145] = 1'b0;
  assign data_mem_pkt_o[146] = 1'b0;
  assign data_mem_pkt_o[147] = 1'b0;
  assign data_mem_pkt_o[148] = 1'b0;
  assign data_mem_pkt_o[149] = 1'b0;
  assign data_mem_pkt_o[150] = 1'b0;
  assign data_mem_pkt_o[151] = 1'b0;
  assign data_mem_pkt_o[152] = 1'b0;
  assign data_mem_pkt_o[153] = 1'b0;
  assign data_mem_pkt_o[154] = 1'b0;
  assign data_mem_pkt_o[155] = 1'b0;
  assign data_mem_pkt_o[156] = 1'b0;
  assign data_mem_pkt_o[157] = 1'b0;
  assign data_mem_pkt_o[158] = 1'b0;
  assign data_mem_pkt_o[159] = 1'b0;
  assign data_mem_pkt_o[160] = 1'b0;
  assign data_mem_pkt_o[161] = 1'b0;
  assign data_mem_pkt_o[162] = 1'b0;
  assign data_mem_pkt_o[163] = 1'b0;
  assign data_mem_pkt_o[164] = 1'b0;
  assign data_mem_pkt_o[165] = 1'b0;
  assign data_mem_pkt_o[166] = 1'b0;
  assign data_mem_pkt_o[167] = 1'b0;
  assign data_mem_pkt_o[168] = 1'b0;
  assign data_mem_pkt_o[169] = 1'b0;
  assign data_mem_pkt_o[170] = 1'b0;
  assign data_mem_pkt_o[171] = 1'b0;
  assign data_mem_pkt_o[172] = 1'b0;
  assign data_mem_pkt_o[173] = 1'b0;
  assign data_mem_pkt_o[174] = 1'b0;
  assign data_mem_pkt_o[175] = 1'b0;
  assign data_mem_pkt_o[176] = 1'b0;
  assign data_mem_pkt_o[177] = 1'b0;
  assign data_mem_pkt_o[178] = 1'b0;
  assign data_mem_pkt_o[179] = 1'b0;
  assign data_mem_pkt_o[180] = 1'b0;
  assign data_mem_pkt_o[181] = 1'b0;
  assign data_mem_pkt_o[182] = 1'b0;
  assign data_mem_pkt_o[183] = 1'b0;
  assign data_mem_pkt_o[184] = 1'b0;
  assign data_mem_pkt_o[185] = 1'b0;
  assign data_mem_pkt_o[186] = 1'b0;
  assign data_mem_pkt_o[187] = 1'b0;
  assign data_mem_pkt_o[188] = 1'b0;
  assign data_mem_pkt_o[189] = 1'b0;
  assign data_mem_pkt_o[190] = 1'b0;
  assign data_mem_pkt_o[191] = 1'b0;
  assign data_mem_pkt_o[192] = 1'b0;
  assign data_mem_pkt_o[193] = 1'b0;
  assign data_mem_pkt_o[194] = 1'b0;
  assign data_mem_pkt_o[195] = 1'b0;
  assign data_mem_pkt_o[196] = 1'b0;
  assign data_mem_pkt_o[197] = 1'b0;
  assign data_mem_pkt_o[198] = 1'b0;
  assign data_mem_pkt_o[199] = 1'b0;
  assign data_mem_pkt_o[200] = 1'b0;
  assign data_mem_pkt_o[201] = 1'b0;
  assign data_mem_pkt_o[202] = 1'b0;
  assign data_mem_pkt_o[203] = 1'b0;
  assign data_mem_pkt_o[204] = 1'b0;
  assign data_mem_pkt_o[205] = 1'b0;
  assign data_mem_pkt_o[206] = 1'b0;
  assign data_mem_pkt_o[207] = 1'b0;
  assign data_mem_pkt_o[208] = 1'b0;
  assign data_mem_pkt_o[209] = 1'b0;
  assign data_mem_pkt_o[210] = 1'b0;
  assign data_mem_pkt_o[211] = 1'b0;
  assign data_mem_pkt_o[212] = 1'b0;
  assign data_mem_pkt_o[213] = 1'b0;
  assign data_mem_pkt_o[214] = 1'b0;
  assign data_mem_pkt_o[215] = 1'b0;
  assign data_mem_pkt_o[216] = 1'b0;
  assign data_mem_pkt_o[217] = 1'b0;
  assign data_mem_pkt_o[218] = 1'b0;
  assign data_mem_pkt_o[219] = 1'b0;
  assign data_mem_pkt_o[220] = 1'b0;
  assign data_mem_pkt_o[221] = 1'b0;
  assign data_mem_pkt_o[222] = 1'b0;
  assign data_mem_pkt_o[223] = 1'b0;
  assign data_mem_pkt_o[224] = 1'b0;
  assign data_mem_pkt_o[225] = 1'b0;
  assign data_mem_pkt_o[226] = 1'b0;
  assign data_mem_pkt_o[227] = 1'b0;
  assign data_mem_pkt_o[228] = 1'b0;
  assign data_mem_pkt_o[229] = 1'b0;
  assign data_mem_pkt_o[230] = 1'b0;
  assign data_mem_pkt_o[231] = 1'b0;
  assign data_mem_pkt_o[232] = 1'b0;
  assign data_mem_pkt_o[233] = 1'b0;
  assign data_mem_pkt_o[234] = 1'b0;
  assign data_mem_pkt_o[235] = 1'b0;
  assign data_mem_pkt_o[236] = 1'b0;
  assign data_mem_pkt_o[237] = 1'b0;
  assign data_mem_pkt_o[238] = 1'b0;
  assign data_mem_pkt_o[239] = 1'b0;
  assign data_mem_pkt_o[240] = 1'b0;
  assign data_mem_pkt_o[241] = 1'b0;
  assign data_mem_pkt_o[242] = 1'b0;
  assign data_mem_pkt_o[243] = 1'b0;
  assign data_mem_pkt_o[244] = 1'b0;
  assign data_mem_pkt_o[245] = 1'b0;
  assign data_mem_pkt_o[246] = 1'b0;
  assign data_mem_pkt_o[247] = 1'b0;
  assign data_mem_pkt_o[248] = 1'b0;
  assign data_mem_pkt_o[249] = 1'b0;
  assign data_mem_pkt_o[250] = 1'b0;
  assign data_mem_pkt_o[251] = 1'b0;
  assign data_mem_pkt_o[252] = 1'b0;
  assign data_mem_pkt_o[253] = 1'b0;
  assign data_mem_pkt_o[254] = 1'b0;
  assign data_mem_pkt_o[255] = 1'b0;
  assign data_mem_pkt_o[256] = 1'b0;
  assign data_mem_pkt_o[257] = 1'b0;
  assign data_mem_pkt_o[258] = 1'b0;
  assign data_mem_pkt_o[259] = 1'b0;
  assign data_mem_pkt_o[260] = 1'b0;
  assign data_mem_pkt_o[261] = 1'b0;
  assign data_mem_pkt_o[262] = 1'b0;
  assign data_mem_pkt_o[263] = 1'b0;
  assign data_mem_pkt_o[264] = 1'b0;
  assign data_mem_pkt_o[265] = 1'b0;
  assign data_mem_pkt_o[266] = 1'b0;
  assign data_mem_pkt_o[267] = 1'b0;
  assign data_mem_pkt_o[268] = 1'b0;
  assign data_mem_pkt_o[269] = 1'b0;
  assign data_mem_pkt_o[270] = 1'b0;
  assign data_mem_pkt_o[271] = 1'b0;
  assign data_mem_pkt_o[272] = 1'b0;
  assign data_mem_pkt_o[273] = 1'b0;
  assign data_mem_pkt_o[274] = 1'b0;
  assign data_mem_pkt_o[275] = 1'b0;
  assign data_mem_pkt_o[276] = 1'b0;
  assign data_mem_pkt_o[277] = 1'b0;
  assign data_mem_pkt_o[278] = 1'b0;
  assign data_mem_pkt_o[279] = 1'b0;
  assign data_mem_pkt_o[280] = 1'b0;
  assign data_mem_pkt_o[281] = 1'b0;
  assign data_mem_pkt_o[282] = 1'b0;
  assign data_mem_pkt_o[283] = 1'b0;
  assign data_mem_pkt_o[284] = 1'b0;
  assign data_mem_pkt_o[285] = 1'b0;
  assign data_mem_pkt_o[286] = 1'b0;
  assign data_mem_pkt_o[287] = 1'b0;
  assign data_mem_pkt_o[288] = 1'b0;
  assign data_mem_pkt_o[289] = 1'b0;
  assign data_mem_pkt_o[290] = 1'b0;
  assign data_mem_pkt_o[291] = 1'b0;
  assign data_mem_pkt_o[292] = 1'b0;
  assign data_mem_pkt_o[293] = 1'b0;
  assign data_mem_pkt_o[294] = 1'b0;
  assign data_mem_pkt_o[295] = 1'b0;
  assign data_mem_pkt_o[296] = 1'b0;
  assign data_mem_pkt_o[297] = 1'b0;
  assign data_mem_pkt_o[298] = 1'b0;
  assign data_mem_pkt_o[299] = 1'b0;
  assign data_mem_pkt_o[300] = 1'b0;
  assign data_mem_pkt_o[301] = 1'b0;
  assign data_mem_pkt_o[302] = 1'b0;
  assign data_mem_pkt_o[303] = 1'b0;
  assign data_mem_pkt_o[304] = 1'b0;
  assign data_mem_pkt_o[305] = 1'b0;
  assign data_mem_pkt_o[306] = 1'b0;
  assign data_mem_pkt_o[307] = 1'b0;
  assign data_mem_pkt_o[308] = 1'b0;
  assign data_mem_pkt_o[309] = 1'b0;
  assign data_mem_pkt_o[310] = 1'b0;
  assign data_mem_pkt_o[311] = 1'b0;
  assign data_mem_pkt_o[312] = 1'b0;
  assign data_mem_pkt_o[313] = 1'b0;
  assign data_mem_pkt_o[314] = 1'b0;
  assign data_mem_pkt_o[315] = 1'b0;
  assign data_mem_pkt_o[316] = 1'b0;
  assign data_mem_pkt_o[317] = 1'b0;
  assign data_mem_pkt_o[318] = 1'b0;
  assign data_mem_pkt_o[319] = 1'b0;
  assign data_mem_pkt_o[320] = 1'b0;
  assign data_mem_pkt_o[321] = 1'b0;
  assign data_mem_pkt_o[322] = 1'b0;
  assign data_mem_pkt_o[323] = 1'b0;
  assign data_mem_pkt_o[324] = 1'b0;
  assign data_mem_pkt_o[325] = 1'b0;
  assign data_mem_pkt_o[326] = 1'b0;
  assign data_mem_pkt_o[327] = 1'b0;
  assign data_mem_pkt_o[328] = 1'b0;
  assign data_mem_pkt_o[329] = 1'b0;
  assign data_mem_pkt_o[330] = 1'b0;
  assign data_mem_pkt_o[331] = 1'b0;
  assign data_mem_pkt_o[332] = 1'b0;
  assign data_mem_pkt_o[333] = 1'b0;
  assign data_mem_pkt_o[334] = 1'b0;
  assign data_mem_pkt_o[335] = 1'b0;
  assign data_mem_pkt_o[336] = 1'b0;
  assign data_mem_pkt_o[337] = 1'b0;
  assign data_mem_pkt_o[338] = 1'b0;
  assign data_mem_pkt_o[339] = 1'b0;
  assign data_mem_pkt_o[340] = 1'b0;
  assign data_mem_pkt_o[341] = 1'b0;
  assign data_mem_pkt_o[342] = 1'b0;
  assign data_mem_pkt_o[343] = 1'b0;
  assign data_mem_pkt_o[344] = 1'b0;
  assign data_mem_pkt_o[345] = 1'b0;
  assign data_mem_pkt_o[346] = 1'b0;
  assign data_mem_pkt_o[347] = 1'b0;
  assign data_mem_pkt_o[348] = 1'b0;
  assign data_mem_pkt_o[349] = 1'b0;
  assign data_mem_pkt_o[350] = 1'b0;
  assign data_mem_pkt_o[351] = 1'b0;
  assign data_mem_pkt_o[352] = 1'b0;
  assign data_mem_pkt_o[353] = 1'b0;
  assign data_mem_pkt_o[354] = 1'b0;
  assign data_mem_pkt_o[355] = 1'b0;
  assign data_mem_pkt_o[356] = 1'b0;
  assign data_mem_pkt_o[357] = 1'b0;
  assign data_mem_pkt_o[358] = 1'b0;
  assign data_mem_pkt_o[359] = 1'b0;
  assign data_mem_pkt_o[360] = 1'b0;
  assign data_mem_pkt_o[361] = 1'b0;
  assign data_mem_pkt_o[362] = 1'b0;
  assign data_mem_pkt_o[363] = 1'b0;
  assign data_mem_pkt_o[364] = 1'b0;
  assign data_mem_pkt_o[365] = 1'b0;
  assign data_mem_pkt_o[366] = 1'b0;
  assign data_mem_pkt_o[367] = 1'b0;
  assign data_mem_pkt_o[368] = 1'b0;
  assign data_mem_pkt_o[369] = 1'b0;
  assign data_mem_pkt_o[370] = 1'b0;
  assign data_mem_pkt_o[371] = 1'b0;
  assign data_mem_pkt_o[372] = 1'b0;
  assign data_mem_pkt_o[373] = 1'b0;
  assign data_mem_pkt_o[374] = 1'b0;
  assign data_mem_pkt_o[375] = 1'b0;
  assign data_mem_pkt_o[376] = 1'b0;
  assign data_mem_pkt_o[377] = 1'b0;
  assign data_mem_pkt_o[378] = 1'b0;
  assign data_mem_pkt_o[379] = 1'b0;
  assign data_mem_pkt_o[380] = 1'b0;
  assign data_mem_pkt_o[381] = 1'b0;
  assign data_mem_pkt_o[382] = 1'b0;
  assign data_mem_pkt_o[383] = 1'b0;
  assign data_mem_pkt_o[384] = 1'b0;
  assign data_mem_pkt_o[385] = 1'b0;
  assign data_mem_pkt_o[386] = 1'b0;
  assign data_mem_pkt_o[387] = 1'b0;
  assign data_mem_pkt_o[388] = 1'b0;
  assign data_mem_pkt_o[389] = 1'b0;
  assign data_mem_pkt_o[390] = 1'b0;
  assign data_mem_pkt_o[391] = 1'b0;
  assign data_mem_pkt_o[392] = 1'b0;
  assign data_mem_pkt_o[393] = 1'b0;
  assign data_mem_pkt_o[394] = 1'b0;
  assign data_mem_pkt_o[395] = 1'b0;
  assign data_mem_pkt_o[396] = 1'b0;
  assign data_mem_pkt_o[397] = 1'b0;
  assign data_mem_pkt_o[398] = 1'b0;
  assign data_mem_pkt_o[399] = 1'b0;
  assign data_mem_pkt_o[400] = 1'b0;
  assign data_mem_pkt_o[401] = 1'b0;
  assign data_mem_pkt_o[402] = 1'b0;
  assign data_mem_pkt_o[403] = 1'b0;
  assign data_mem_pkt_o[404] = 1'b0;
  assign data_mem_pkt_o[405] = 1'b0;
  assign data_mem_pkt_o[406] = 1'b0;
  assign data_mem_pkt_o[407] = 1'b0;
  assign data_mem_pkt_o[408] = 1'b0;
  assign data_mem_pkt_o[409] = 1'b0;
  assign data_mem_pkt_o[410] = 1'b0;
  assign data_mem_pkt_o[411] = 1'b0;
  assign data_mem_pkt_o[412] = 1'b0;
  assign data_mem_pkt_o[413] = 1'b0;
  assign data_mem_pkt_o[414] = 1'b0;
  assign data_mem_pkt_o[415] = 1'b0;
  assign data_mem_pkt_o[416] = 1'b0;
  assign data_mem_pkt_o[417] = 1'b0;
  assign data_mem_pkt_o[418] = 1'b0;
  assign data_mem_pkt_o[419] = 1'b0;
  assign data_mem_pkt_o[420] = 1'b0;
  assign data_mem_pkt_o[421] = 1'b0;
  assign data_mem_pkt_o[422] = 1'b0;
  assign data_mem_pkt_o[423] = 1'b0;
  assign data_mem_pkt_o[424] = 1'b0;
  assign data_mem_pkt_o[425] = 1'b0;
  assign data_mem_pkt_o[426] = 1'b0;
  assign data_mem_pkt_o[427] = 1'b0;
  assign data_mem_pkt_o[428] = 1'b0;
  assign data_mem_pkt_o[429] = 1'b0;
  assign data_mem_pkt_o[430] = 1'b0;
  assign data_mem_pkt_o[431] = 1'b0;
  assign data_mem_pkt_o[432] = 1'b0;
  assign data_mem_pkt_o[433] = 1'b0;
  assign data_mem_pkt_o[434] = 1'b0;
  assign data_mem_pkt_o[435] = 1'b0;
  assign data_mem_pkt_o[436] = 1'b0;
  assign data_mem_pkt_o[437] = 1'b0;
  assign data_mem_pkt_o[438] = 1'b0;
  assign data_mem_pkt_o[439] = 1'b0;
  assign data_mem_pkt_o[440] = 1'b0;
  assign data_mem_pkt_o[441] = 1'b0;
  assign data_mem_pkt_o[442] = 1'b0;
  assign data_mem_pkt_o[443] = 1'b0;
  assign data_mem_pkt_o[444] = 1'b0;
  assign data_mem_pkt_o[445] = 1'b0;
  assign data_mem_pkt_o[446] = 1'b0;
  assign data_mem_pkt_o[447] = 1'b0;
  assign data_mem_pkt_o[448] = 1'b0;
  assign data_mem_pkt_o[449] = 1'b0;
  assign data_mem_pkt_o[450] = 1'b0;
  assign data_mem_pkt_o[451] = 1'b0;
  assign data_mem_pkt_o[452] = 1'b0;
  assign data_mem_pkt_o[453] = 1'b0;
  assign data_mem_pkt_o[454] = 1'b0;
  assign data_mem_pkt_o[455] = 1'b0;
  assign data_mem_pkt_o[456] = 1'b0;
  assign data_mem_pkt_o[457] = 1'b0;
  assign data_mem_pkt_o[458] = 1'b0;
  assign data_mem_pkt_o[459] = 1'b0;
  assign data_mem_pkt_o[460] = 1'b0;
  assign data_mem_pkt_o[461] = 1'b0;
  assign data_mem_pkt_o[462] = 1'b0;
  assign data_mem_pkt_o[463] = 1'b0;
  assign data_mem_pkt_o[464] = 1'b0;
  assign data_mem_pkt_o[465] = 1'b0;
  assign data_mem_pkt_o[466] = 1'b0;
  assign data_mem_pkt_o[467] = 1'b0;
  assign data_mem_pkt_o[468] = 1'b0;
  assign data_mem_pkt_o[469] = 1'b0;
  assign data_mem_pkt_o[470] = 1'b0;
  assign data_mem_pkt_o[471] = 1'b0;
  assign data_mem_pkt_o[472] = 1'b0;
  assign data_mem_pkt_o[473] = 1'b0;
  assign data_mem_pkt_o[474] = 1'b0;
  assign data_mem_pkt_o[475] = 1'b0;
  assign data_mem_pkt_o[476] = 1'b0;
  assign data_mem_pkt_o[477] = 1'b0;
  assign data_mem_pkt_o[478] = 1'b0;
  assign data_mem_pkt_o[479] = 1'b0;
  assign data_mem_pkt_o[480] = 1'b0;
  assign data_mem_pkt_o[481] = 1'b0;
  assign data_mem_pkt_o[482] = 1'b0;
  assign data_mem_pkt_o[483] = 1'b0;
  assign data_mem_pkt_o[484] = 1'b0;
  assign data_mem_pkt_o[485] = 1'b0;
  assign data_mem_pkt_o[486] = 1'b0;
  assign data_mem_pkt_o[487] = 1'b0;
  assign data_mem_pkt_o[488] = 1'b0;
  assign data_mem_pkt_o[489] = 1'b0;
  assign data_mem_pkt_o[490] = 1'b0;
  assign data_mem_pkt_o[491] = 1'b0;
  assign data_mem_pkt_o[492] = 1'b0;
  assign data_mem_pkt_o[493] = 1'b0;
  assign data_mem_pkt_o[494] = 1'b0;
  assign data_mem_pkt_o[495] = 1'b0;
  assign data_mem_pkt_o[496] = 1'b0;
  assign data_mem_pkt_o[497] = 1'b0;
  assign data_mem_pkt_o[498] = 1'b0;
  assign data_mem_pkt_o[499] = 1'b0;
  assign data_mem_pkt_o[500] = 1'b0;
  assign data_mem_pkt_o[501] = 1'b0;
  assign data_mem_pkt_o[502] = 1'b0;
  assign data_mem_pkt_o[503] = 1'b0;
  assign data_mem_pkt_o[504] = 1'b0;
  assign data_mem_pkt_o[505] = 1'b0;
  assign data_mem_pkt_o[506] = 1'b0;
  assign data_mem_pkt_o[507] = 1'b0;
  assign data_mem_pkt_o[508] = 1'b0;
  assign data_mem_pkt_o[509] = 1'b0;
  assign data_mem_pkt_o[510] = 1'b0;
  assign data_mem_pkt_o[511] = 1'b0;
  assign data_mem_pkt_o[512] = 1'b0;
  assign lce_resp_o[23] = 1'b0;
  assign lce_tr_resp_o[537] = lce_id_i[0];
  assign lce_data_resp_o[535] = lce_id_i[0];
  assign lce_resp_o[24] = lce_id_i[0];
  assign N31 = N28 & N29;
  assign N32 = N31 & N30;
  assign N33 = state_r[2] | state_r[1];
  assign N34 = N33 | N30;
  assign N36 = state_r[2] | N29;
  assign N37 = N36 | state_r[0];
  assign N39 = state_r[2] | N29;
  assign N40 = N39 | N30;
  assign N42 = N28 | state_r[1];
  assign N43 = N42 | state_r[0];
  assign N45 = N28 | state_r[1];
  assign N46 = N45 | N30;
  assign N48 = state_r[2] & state_r[1];
  assign N49 = N86 & N75;
  assign N50 = lce_cmd_i[33] | lce_cmd_i[32];
  assign N51 = N50 | N75;
  assign N68 = N70 | lce_cmd_i[31];
  assign N70 = lce_cmd_i[33] | N80;
  assign N71 = N70 | N75;
  assign N73 = N76 | lce_cmd_i[31];
  assign N76 = N79 | lce_cmd_i[32];
  assign N77 = N76 | N75;
  assign N81 = N79 | N80;
  assign N82 = N81 | lce_cmd_i[31];
  assign N84 = lce_cmd_i[33] & lce_cmd_i[32];
  assign N85 = N84 & lce_cmd_i[31];
  assign N86 = N79 & N80;
  assign N698 = (N690)? dirty_i[0] : 
                (N692)? dirty_i[1] : 
                (N694)? dirty_i[2] : 
                (N696)? dirty_i[3] : 
                (N691)? dirty_i[4] : 
                (N693)? dirty_i[5] : 
                (N695)? dirty_i[6] : 
                (N697)? dirty_i[7] : 1'b0;
  assign N1604 = state_r[1] | state_r[2];
  assign lce_sync_done_o = state_r[0] | N1604;
  assign N1606 = ~sync_ack_count_r[0];
  assign N55 = sync_ack_count_r[0] ^ 1'b1;
  assign N58 = (N0)? lce_cmd_i[34] : 
               (N1)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N0 = N49;
  assign N1 = N52;
  assign N2 = N53;
  assign N59 = (N0)? lce_cmd_v_i : 
               (N1)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N60 = (N0)? lce_resp_yumi_i : 
               (N1)? N57 : 
               (N2)? 1'b0 : 1'b0;
  assign { N66, N65, N64, N63, N62, N61 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N1)? lce_cmd_i[20:15] : 
                                            (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N67 = (N0)? 1'b0 : 
               (N1)? lce_cmd_v_i : 
               (N2)? 1'b0 : 1'b0;
  assign N90 = (N3)? 1'b0 : 
               (N4)? lce_cmd_v_i : 1'b0;
  assign N3 = invalidated_tag_r;
  assign N4 = N89;
  assign N93 = (N5)? 1'b0 : 
               (N1237)? 1'b1 : 
               (N92)? tag_mem_pkt_yumi_i : 1'b0;
  assign N5 = lce_resp_yumi_i;
  assign { N103, N102, N101, N100, N99, N98, N97, N96, N95 } = (N6)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                                               (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = N69;
  assign N7 = N72;
  assign N8 = N74;
  assign N9 = N78;
  assign N10 = N83;
  assign N11 = N87;
  assign N104 = (N6)? lce_cmd_v_i : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 1'b0;
  assign { N106, N105 } = (N6)? { data_mem_pkt_yumi_i, N88 } : 
                          (N7)? { stat_mem_pkt_yumi_i, 1'b1 } : 1'b0;
  assign { N116, N115, N114, N113, N112, N111, N110, N109, N108, N107 } = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N7)? { lce_cmd_i[20:15], lce_cmd_i[8:6], 1'b1 } : 
                                                                          (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N117 = (N6)? 1'b0 : 
                (N7)? lce_cmd_v_i : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 1'b0;
  assign { N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118 } = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                  (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                  (N8)? { lce_cmd_i[20:15], lce_cmd_i[8:4], lce_cmd_i[30:21], 1'b1 } : 
                                                                                                                                                  (N9)? { lce_cmd_i[20:15], lce_cmd_i[8:4], lce_cmd_i[30:21], 1'b1 } : 
                                                                                                                                                  (N10)? { lce_cmd_i[20:15], lce_cmd_i[8:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                  (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N140 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? lce_cmd_v_i : 
                (N9)? lce_cmd_v_i : 
                (N10)? N90 : 
                (N11)? 1'b0 : 1'b0;
  assign N141 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? tag_mem_pkt_yumi_i : 
                (N9)? tag_mem_pkt_yumi_i : 
                (N10)? lce_resp_yumi_i : 
                (N11)? 1'b0 : 1'b0;
  assign N142 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? tag_mem_pkt_yumi_i : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 1'b0;
  assign N143 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? tag_mem_pkt_yumi_i : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 1'b0;
  assign { N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144 } = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                              (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                              (N10)? { lce_cmd_i[34:34], 1'b1, lce_cmd_i[30:9] } : 
                                                                                                                                                              (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N168 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? N94 : 
                (N11)? 1'b0 : 1'b0;
  assign { N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171 } = (N12)? data_buf_r : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N13)? data_mem_data_i : 1'b0;
  assign N12 = tr_data_buffered_r;
  assign N13 = N170;
  assign N699 = ~N698;
  assign N710 = (N14)? 1'b0 : 
                (N1241)? 1'b1 : 
                (N709)? wb_data_read_r : 1'b0;
  assign N14 = lce_data_resp_done;
  assign N713 = (N14)? 1'b0 : 
                (N1242)? 1'b1 : 
                (N712)? data_mem_pkt_yumi_i : 1'b0;
  assign N716 = (N15)? 1'b0 : 
                (N16)? N715 : 1'b0;
  assign N15 = wb_dirty_cleared_r;
  assign N16 = N714;
  assign N719 = (N14)? 1'b0 : 
                (N1243)? 1'b1 : 
                (N718)? stat_mem_pkt_yumi_i : 1'b0;
  assign { N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721 } = (N17)? data_buf_r : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       (N18)? data_mem_data_i : 1'b0;
  assign N17 = wb_data_buffered_r;
  assign N18 = N720;
  assign stat_mem_pkt_o[0] = (N19)? N107 : 
                             (N1235)? 1'b0 : 1'b0;
  assign N19 = N35;
  assign stat_mem_pkt_o[10:2] = (N20)? { N66, N65, N64, N63, N62, N61, 1'b0, 1'b0, 1'b0 } : 
                                (N19)? { N116, N115, N114, N113, N112, N111, N110, N109, N108 } : 
                                (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                (N23)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = N32;
  assign N21 = N38;
  assign N22 = N41;
  assign N23 = stat_mem_pkt_o[1];
  assign N24 = N47;
  assign N25 = N48;
  assign stat_mem_pkt_v_o = (N20)? N67 : 
                            (N19)? N117 : 
                            (N21)? 1'b0 : 
                            (N22)? 1'b0 : 
                            (N23)? N716 : 
                            (N24)? 1'b0 : 
                            (N25)? 1'b0 : 1'b0;
  assign { lce_resp_o[25:25], lce_resp_o[22:0] } = (N20)? { N58, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N19)? { N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144 } : 
                                                   (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_resp_v_o = (N20)? N59 : 
                        (N19)? N168 : 
                        (N21)? 1'b0 : 
                        (N22)? 1'b0 : 
                        (N23)? 1'b0 : 
                        (N24)? 1'b0 : 
                        (N25)? 1'b0 : 1'b0;
  assign lce_cmd_yumi_o = (N20)? N60 : 
                          (N19)? N141 : 
                          (N21)? lce_tr_resp_done : 
                          (N22)? 1'b0 : 
                          (N23)? lce_data_resp_done : 
                          (N24)? lce_data_resp_done : 
                          (N25)? 1'b0 : 1'b0;
  assign state_n = (N20)? { 1'b0, 1'b0, N56 } : 
                   (N19)? { 1'b0, N106, N105 } : 
                   (N21)? { 1'b0, N169, lce_tr_resp_done } : 
                   (N22)? { 1'b1, 1'b0, N699 } : 
                   (N23)? { N1234, 1'b0, lce_data_resp_done } : 
                   (N24)? { N1234, 1'b0, 1'b1 } : 
                   (N25)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_pkt_o = (N20)? { N66, N65, N64, N63, N62, N61, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N19)? { N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N83 } : 
                         (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_pkt_v_o = (N20)? N67 : 
                           (N19)? N140 : 
                           (N21)? 1'b0 : 
                           (N22)? 1'b0 : 
                           (N23)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N25)? 1'b0 : 1'b0;
  assign data_mem_pkt_o[521:513] = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N19)? { N103, N102, N101, N100, N99, N98, N97, N96, N95 } : 
                                   (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N23)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                   (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign data_mem_pkt_v_o = (N20)? 1'b0 : 
                            (N19)? N104 : 
                            (N21)? 1'b0 : 
                            (N22)? 1'b0 : 
                            (N23)? N700 : 
                            (N24)? 1'b0 : 
                            (N25)? 1'b0 : 1'b0;
  assign tag_set_o = (N20)? 1'b0 : 
                     (N19)? N142 : 
                     (N21)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N25)? 1'b0 : 1'b0;
  assign tag_set_wakeup_o = (N20)? 1'b0 : 
                            (N19)? N143 : 
                            (N21)? 1'b0 : 
                            (N22)? 1'b0 : 
                            (N23)? 1'b0 : 
                            (N24)? 1'b0 : 
                            (N25)? 1'b0 : 1'b0;
  assign { lce_tr_resp_o[538:538], lce_tr_resp_o[536:0] } = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N21)? { lce_cmd_i[3:0], lce_cmd_i[30:9], N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171 } : 
                                                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_tr_resp_v_o = (N20)? 1'b0 : 
                           (N19)? 1'b0 : 
                           (N21)? 1'b1 : 
                           (N22)? 1'b0 : 
                           (N23)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N25)? 1'b0 : 1'b0;
  assign { lce_data_resp_o[536:536], lce_data_resp_o[534:0] } = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N23)? { lce_cmd_i[34:34], 1'b0, lce_cmd_i[30:9], N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721 } : 
                                                                (N24)? { lce_cmd_i[34:34], 1'b1, lce_cmd_i[30:9], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_data_resp_v_o = (N20)? 1'b0 : 
                             (N19)? 1'b0 : 
                             (N21)? 1'b0 : 
                             (N22)? 1'b0 : 
                             (N23)? N1233 : 
                             (N24)? 1'b1 : 
                             (N25)? 1'b0 : 1'b0;
  assign { N1247, N1246, N1245 } = (N26)? { 1'b0, 1'b0, 1'b0 } : 
                                   (N27)? state_n : 1'b0;
  assign N26 = reset_i;
  assign N27 = N1244;
  assign N1248 = (N26)? 1'b0 : 
                 (N27)? N55 : 1'b0;
  assign N1249 = (N26)? 1'b0 : 
                 (N27)? N169 : 1'b0;
  assign N1250 = (N26)? 1'b0 : 
                 (N27)? N710 : 1'b0;
  assign N1251 = (N26)? 1'b0 : 
                 (N27)? N713 : 1'b0;
  assign N1252 = (N26)? 1'b0 : 
                 (N27)? N719 : 1'b0;
  assign N1253 = (N26)? 1'b0 : 
                 (N27)? N93 : 1'b0;
  assign lce_tr_resp_done = lce_tr_resp_v_o & lce_tr_resp_ready_i;
  assign lce_data_resp_done = lce_data_resp_ready_i & lce_data_resp_v_o;
  assign N28 = ~state_r[2];
  assign N29 = ~state_r[1];
  assign N30 = ~state_r[0];
  assign N35 = ~N34;
  assign N38 = ~N37;
  assign N41 = ~N40;
  assign N44 = ~N43;
  assign N47 = ~N46;
  assign stat_mem_pkt_o[1] = N44;
  assign N52 = ~N51;
  assign N53 = lce_cmd_i[33] | lce_cmd_i[32];
  assign N54 = ~lce_resp_yumi_i;
  assign N56 = N1606 & lce_resp_yumi_i;
  assign N57 = tag_mem_pkt_yumi_i & stat_mem_pkt_yumi_i;
  assign N69 = ~N68;
  assign N72 = ~N71;
  assign N74 = ~N73;
  assign N75 = ~lce_cmd_i[31];
  assign N78 = ~N77;
  assign N79 = ~lce_cmd_i[33];
  assign N80 = ~lce_cmd_i[32];
  assign N83 = ~N82;
  assign N87 = N85 | N86;
  assign N88 = ~data_mem_pkt_yumi_i;
  assign N89 = ~invalidated_tag_r;
  assign N91 = invalidated_tag_r | lce_resp_yumi_i;
  assign N92 = ~N91;
  assign N94 = invalidated_tag_r | tag_mem_pkt_yumi_i;
  assign N169 = ~lce_tr_resp_done;
  assign N170 = ~tr_data_buffered_r;
  assign N683 = ~lce_cmd_i[6];
  assign N684 = ~lce_cmd_i[7];
  assign N685 = N683 & N684;
  assign N686 = N683 & lce_cmd_i[7];
  assign N687 = lce_cmd_i[6] & N684;
  assign N688 = lce_cmd_i[6] & lce_cmd_i[7];
  assign N689 = ~lce_cmd_i[8];
  assign N690 = N685 & N689;
  assign N691 = N685 & lce_cmd_i[8];
  assign N692 = N687 & N689;
  assign N693 = N687 & lce_cmd_i[8];
  assign N694 = N686 & N689;
  assign N695 = N686 & lce_cmd_i[8];
  assign N696 = N688 & N689;
  assign N697 = N688 & lce_cmd_i[8];
  assign N700 = ~wb_data_read_r;
  assign N701 = ~N1239;
  assign N702 = N701;
  assign N703 = N701;
  assign N704 = N701;
  assign N705 = N701;
  assign N706 = N701;
  assign N707 = N701;
  assign N708 = wb_data_buffered_r | lce_data_resp_done;
  assign N709 = ~N708;
  assign N711 = wb_data_read_r | lce_data_resp_done;
  assign N712 = ~N711;
  assign N714 = ~wb_dirty_cleared_r;
  assign N715 = wb_data_read_r | data_mem_pkt_yumi_i;
  assign N717 = wb_dirty_cleared_r | lce_data_resp_done;
  assign N718 = ~N717;
  assign N720 = ~wb_data_buffered_r;
  assign N1233 = wb_data_read_r & N1607;
  assign N1607 = wb_dirty_cleared_r | stat_mem_pkt_yumi_i;
  assign N1234 = ~lce_data_resp_done;
  assign N1235 = N34;
  assign N1236 = ~lce_resp_yumi_i;
  assign N1237 = invalidated_tag_r & N1236;
  assign N1238 = ~wb_data_buffered_r;
  assign N1239 = wb_data_read_r & N1238;
  assign N1240 = ~lce_data_resp_done;
  assign N1241 = wb_data_buffered_r & N1240;
  assign N1242 = wb_data_read_r & N1240;
  assign N1243 = wb_dirty_cleared_r & N1240;
  assign N1244 = ~reset_i;
  assign N1254 = N32 & N1244;
  assign N1255 = N35 & N1244;
  assign N1256 = N1254 | N1255;
  assign N1257 = N38 & N1244;
  assign N1258 = tr_data_buffered_r & N1257;
  assign N1259 = N1256 | N1258;
  assign N1260 = N41 & N1244;
  assign N1261 = N1259 | N1260;
  assign N1262 = stat_mem_pkt_o[1] & N1244;
  assign N1263 = N702 & N1262;
  assign N1264 = N1261 | N1263;
  assign N1265 = N47 & N1244;
  assign N1266 = N1264 | N1265;
  assign N1267 = N48 & N1244;
  assign N1268 = N1266 | N1267;
  assign N1269 = ~N1268;
  assign N1270 = N1244 & N1269;
  assign N1271 = N32 & N1244;
  assign N1272 = N35 & N1244;
  assign N1273 = N1271 | N1272;
  assign N1274 = N38 & N1244;
  assign N1275 = tr_data_buffered_r & N1274;
  assign N1276 = N1273 | N1275;
  assign N1277 = N41 & N1244;
  assign N1278 = N1276 | N1277;
  assign N1279 = stat_mem_pkt_o[1] & N1244;
  assign N1280 = N702 & N1279;
  assign N1281 = N1278 | N1280;
  assign N1282 = N47 & N1244;
  assign N1283 = N1281 | N1282;
  assign N1284 = N48 & N1244;
  assign N1285 = N1283 | N1284;
  assign N1286 = ~N1285;
  assign N1287 = N1244 & N1286;
  assign N1288 = N32 & N1244;
  assign N1289 = N35 & N1244;
  assign N1290 = N1288 | N1289;
  assign N1291 = N38 & N1244;
  assign N1292 = tr_data_buffered_r & N1291;
  assign N1293 = N1290 | N1292;
  assign N1294 = N41 & N1244;
  assign N1295 = N1293 | N1294;
  assign N1296 = stat_mem_pkt_o[1] & N1244;
  assign N1297 = N702 & N1296;
  assign N1298 = N1295 | N1297;
  assign N1299 = N47 & N1244;
  assign N1300 = N1298 | N1299;
  assign N1301 = N48 & N1244;
  assign N1302 = N1300 | N1301;
  assign N1303 = ~N1302;
  assign N1304 = N1244 & N1303;
  assign N1305 = N32 & N1244;
  assign N1306 = N35 & N1244;
  assign N1307 = N1305 | N1306;
  assign N1308 = N38 & N1244;
  assign N1309 = tr_data_buffered_r & N1308;
  assign N1310 = N1307 | N1309;
  assign N1311 = N41 & N1244;
  assign N1312 = N1310 | N1311;
  assign N1313 = stat_mem_pkt_o[1] & N1244;
  assign N1314 = N702 & N1313;
  assign N1315 = N1312 | N1314;
  assign N1316 = N47 & N1244;
  assign N1317 = N1315 | N1316;
  assign N1318 = N48 & N1244;
  assign N1319 = N1317 | N1318;
  assign N1320 = ~N1319;
  assign N1321 = N1244 & N1320;
  assign N1322 = N32 & N1244;
  assign N1323 = N35 & N1244;
  assign N1324 = N1322 | N1323;
  assign N1325 = N38 & N1244;
  assign N1326 = tr_data_buffered_r & N1325;
  assign N1327 = N1324 | N1326;
  assign N1328 = N41 & N1244;
  assign N1329 = N1327 | N1328;
  assign N1330 = stat_mem_pkt_o[1] & N1244;
  assign N1331 = N702 & N1330;
  assign N1332 = N1329 | N1331;
  assign N1333 = N47 & N1244;
  assign N1334 = N1332 | N1333;
  assign N1335 = N48 & N1244;
  assign N1336 = N1334 | N1335;
  assign N1337 = ~N1336;
  assign N1338 = N1244 & N1337;
  assign N1339 = N32 & N1244;
  assign N1340 = N35 & N1244;
  assign N1341 = N1339 | N1340;
  assign N1342 = N38 & N1244;
  assign N1343 = tr_data_buffered_r & N1342;
  assign N1344 = N1341 | N1343;
  assign N1345 = N41 & N1244;
  assign N1346 = N1344 | N1345;
  assign N1347 = stat_mem_pkt_o[1] & N1244;
  assign N1348 = N702 & N1347;
  assign N1349 = N1346 | N1348;
  assign N1350 = N47 & N1244;
  assign N1351 = N1349 | N1350;
  assign N1352 = N48 & N1244;
  assign N1353 = N1351 | N1352;
  assign N1354 = ~N1353;
  assign N1355 = N1244 & N1354;
  assign N1356 = N1346 | N1331;
  assign N1357 = N1356 | N1350;
  assign N1358 = N1357 | N1352;
  assign N1359 = ~N1358;
  assign N1360 = N1244 & N1359;
  assign N1361 = N1341 | N1326;
  assign N1362 = N1361 | N1345;
  assign N1363 = N1362 | N1331;
  assign N1364 = N1363 | N1350;
  assign N1365 = N1364 | N1352;
  assign N1366 = ~N1365;
  assign N1367 = N1244 & N1366;
  assign N1368 = N1361 | N1328;
  assign N1369 = N1368 | N1331;
  assign N1370 = N1369 | N1333;
  assign N1371 = N1370 | N1335;
  assign N1372 = ~N1371;
  assign N1373 = N1244 & N1372;
  assign N1374 = N1322 | N1340;
  assign N1375 = N1374 | N1326;
  assign N1376 = N1375 | N1328;
  assign N1377 = N1376 | N1331;
  assign N1378 = N1377 | N1333;
  assign N1379 = N1378 | N1335;
  assign N1380 = ~N1379;
  assign N1381 = N1244 & N1380;
  assign N1382 = N703 & N1330;
  assign N1383 = N1329 | N1382;
  assign N1384 = N1383 | N1333;
  assign N1385 = N1384 | N1335;
  assign N1386 = ~N1385;
  assign N1387 = N1244 & N1386;
  assign N1388 = N703 & N1313;
  assign N1389 = N1329 | N1388;
  assign N1390 = N1389 | N1333;
  assign N1391 = N1390 | N1335;
  assign N1392 = ~N1391;
  assign N1393 = N1244 & N1392;
  assign N1394 = N1324 | N1309;
  assign N1395 = N1394 | N1328;
  assign N1396 = N1395 | N1388;
  assign N1397 = N1396 | N1333;
  assign N1398 = N1397 | N1335;
  assign N1399 = ~N1398;
  assign N1400 = N1244 & N1399;
  assign N1401 = N1394 | N1311;
  assign N1402 = N1401 | N1388;
  assign N1403 = N1402 | N1316;
  assign N1404 = N1403 | N1318;
  assign N1405 = ~N1404;
  assign N1406 = N1244 & N1405;
  assign N1407 = N1305 | N1323;
  assign N1408 = N1407 | N1309;
  assign N1409 = N1408 | N1311;
  assign N1410 = N1409 | N1388;
  assign N1411 = N1410 | N1316;
  assign N1412 = N1411 | N1318;
  assign N1413 = ~N1412;
  assign N1414 = N1244 & N1413;
  assign N1415 = N1312 | N1388;
  assign N1416 = N1415 | N1316;
  assign N1417 = N1416 | N1318;
  assign N1418 = ~N1417;
  assign N1419 = N1244 & N1418;
  assign N1420 = N704 & N1313;
  assign N1421 = N1312 | N1420;
  assign N1422 = N1421 | N1316;
  assign N1423 = N1422 | N1318;
  assign N1424 = ~N1423;
  assign N1425 = N1244 & N1424;
  assign N1426 = N704 & N1296;
  assign N1427 = N1312 | N1426;
  assign N1428 = N1427 | N1316;
  assign N1429 = N1428 | N1318;
  assign N1430 = ~N1429;
  assign N1431 = N1244 & N1430;
  assign N1432 = N1307 | N1292;
  assign N1433 = N1432 | N1311;
  assign N1434 = N1433 | N1426;
  assign N1435 = N1434 | N1316;
  assign N1436 = N1435 | N1318;
  assign N1437 = ~N1436;
  assign N1438 = N1244 & N1437;
  assign N1439 = N1432 | N1294;
  assign N1440 = N1439 | N1426;
  assign N1441 = N1440 | N1299;
  assign N1442 = N1441 | N1301;
  assign N1443 = ~N1442;
  assign N1444 = N1244 & N1443;
  assign N1445 = N1288 | N1306;
  assign N1446 = N1445 | N1292;
  assign N1447 = N1446 | N1294;
  assign N1448 = N1447 | N1426;
  assign N1449 = N1448 | N1299;
  assign N1450 = N1449 | N1301;
  assign N1451 = ~N1450;
  assign N1452 = N1244 & N1451;
  assign N1453 = N1295 | N1426;
  assign N1454 = N1453 | N1299;
  assign N1455 = N1454 | N1301;
  assign N1456 = ~N1455;
  assign N1457 = N1244 & N1456;
  assign N1458 = N705 & N1296;
  assign N1459 = N1295 | N1458;
  assign N1460 = N1459 | N1299;
  assign N1461 = N1460 | N1301;
  assign N1462 = ~N1461;
  assign N1463 = N1244 & N1462;
  assign N1464 = N705 & N1279;
  assign N1465 = N1295 | N1464;
  assign N1466 = N1465 | N1299;
  assign N1467 = N1466 | N1301;
  assign N1468 = ~N1467;
  assign N1469 = N1244 & N1468;
  assign N1470 = N1290 | N1275;
  assign N1471 = N1470 | N1294;
  assign N1472 = N1471 | N1464;
  assign N1473 = N1472 | N1299;
  assign N1474 = N1473 | N1301;
  assign N1475 = ~N1474;
  assign N1476 = N1244 & N1475;
  assign N1477 = N1470 | N1277;
  assign N1478 = N1477 | N1464;
  assign N1479 = N1478 | N1282;
  assign N1480 = N1479 | N1284;
  assign N1481 = ~N1480;
  assign N1482 = N1244 & N1481;
  assign N1483 = N1271 | N1289;
  assign N1484 = N1483 | N1275;
  assign N1485 = N1484 | N1277;
  assign N1486 = N1485 | N1464;
  assign N1487 = N1486 | N1282;
  assign N1488 = N1487 | N1284;
  assign N1489 = ~N1488;
  assign N1490 = N1244 & N1489;
  assign N1491 = N1278 | N1464;
  assign N1492 = N1491 | N1282;
  assign N1493 = N1492 | N1284;
  assign N1494 = ~N1493;
  assign N1495 = N1244 & N1494;
  assign N1496 = N706 & N1279;
  assign N1497 = N1278 | N1496;
  assign N1498 = N1497 | N1282;
  assign N1499 = N1498 | N1284;
  assign N1500 = ~N1499;
  assign N1501 = N1244 & N1500;
  assign N1502 = N706 & N1262;
  assign N1503 = N1278 | N1502;
  assign N1504 = N1503 | N1282;
  assign N1505 = N1504 | N1284;
  assign N1506 = ~N1505;
  assign N1507 = N1244 & N1506;
  assign N1508 = N1273 | N1258;
  assign N1509 = N1508 | N1277;
  assign N1510 = N1509 | N1502;
  assign N1511 = N1510 | N1282;
  assign N1512 = N1511 | N1284;
  assign N1513 = ~N1512;
  assign N1514 = N1244 & N1513;
  assign N1515 = N1508 | N1260;
  assign N1516 = N1515 | N1502;
  assign N1517 = N1516 | N1265;
  assign N1518 = N1517 | N1267;
  assign N1519 = ~N1518;
  assign N1520 = N1244 & N1519;
  assign N1521 = N1254 | N1272;
  assign N1522 = N1521 | N1258;
  assign N1523 = N1522 | N1260;
  assign N1524 = N1523 | N1502;
  assign N1525 = N1524 | N1265;
  assign N1526 = N1525 | N1267;
  assign N1527 = ~N1526;
  assign N1528 = N1244 & N1527;
  assign N1529 = N1261 | N1502;
  assign N1530 = N1529 | N1265;
  assign N1531 = N1530 | N1267;
  assign N1532 = ~N1531;
  assign N1533 = N1244 & N1532;
  assign N1534 = N707 & N1262;
  assign N1535 = N1261 | N1534;
  assign N1536 = N1535 | N1265;
  assign N1537 = N1536 | N1267;
  assign N1538 = ~N1537;
  assign N1539 = N1244 & N1538;
  assign N1540 = N705 & N1262;
  assign N1541 = N1261 | N1540;
  assign N1542 = N1541 | N1265;
  assign N1543 = N1542 | N1267;
  assign N1544 = ~N1543;
  assign N1545 = N1244 & N1544;
  assign N1546 = N704 & N1262;
  assign N1547 = N1261 | N1546;
  assign N1548 = N1547 | N1265;
  assign N1549 = N1548 | N1267;
  assign N1550 = ~N1549;
  assign N1551 = N1244 & N1550;
  assign N1552 = N703 & N1262;
  assign N1553 = N1261 | N1552;
  assign N1554 = N1553 | N1265;
  assign N1555 = N1554 | N1267;
  assign N1556 = ~N1555;
  assign N1557 = N1244 & N1556;
  assign N1558 = N52 & N1254;
  assign N1559 = N53 & N1254;
  assign N1560 = N1558 | N1559;
  assign N1561 = N74 & N1255;
  assign N1562 = N1560 | N1561;
  assign N1563 = N78 & N1255;
  assign N1564 = N1562 | N1563;
  assign N1565 = N83 & N1255;
  assign N1566 = N1564 | N1565;
  assign N1567 = N87 & N1255;
  assign N1568 = N1566 | N1567;
  assign N1569 = ~N1568;
  assign N1570 = N49 & N1254;
  assign N1571 = N54 & N1570;
  assign N1572 = N1571 | N1558;
  assign N1573 = N1572 | N1559;
  assign N1574 = N1573 | N1255;
  assign N1575 = N1574 | N1257;
  assign N1576 = N1575 | N1260;
  assign N1577 = N1576 | N1262;
  assign N1578 = N1577 | N1265;
  assign N1579 = N1578 | N1267;
  assign N1580 = ~N1579;
  assign N1581 = N1256 | N1260;
  assign N1582 = N1581 | N1262;
  assign N1583 = N1582 | N1265;
  assign N1584 = N1583 | N1267;
  assign N1585 = ~N1584;
  assign N1586 = N1256 | N1257;
  assign N1587 = N1586 | N1260;
  assign N1588 = N1587 | N1265;
  assign N1589 = N1588 | N1267;
  assign N1590 = ~N1589;
  assign N1591 = N69 & N1255;
  assign N1592 = N1254 | N1591;
  assign N1593 = N72 & N1255;
  assign N1594 = N1592 | N1593;
  assign N1595 = N1594 | N1561;
  assign N1596 = N1595 | N1563;
  assign N1597 = N1596 | N1567;
  assign N1598 = N1597 | N1257;
  assign N1599 = N1598 | N1260;
  assign N1600 = N1599 | N1262;
  assign N1601 = N1600 | N1265;
  assign N1602 = N1601 | N1267;
  assign N1603 = ~N1602;

  always @(posedge clk_i) begin
    if(N1270) begin
      { data_buf_r[511:511], data_buf_r[0:0] } <= { data_mem_data_i[511:511], data_mem_data_i[0:0] };
    end 
    if(N1287) begin
      { data_buf_r[510:510] } <= { data_mem_data_i[510:510] };
    end 
    if(N1304) begin
      { data_buf_r[509:509] } <= { data_mem_data_i[509:509] };
    end 
    if(N1321) begin
      { data_buf_r[508:508] } <= { data_mem_data_i[508:508] };
    end 
    if(N1338) begin
      { data_buf_r[507:507], data_buf_r[472:413] } <= { data_mem_data_i[507:507], data_mem_data_i[472:413] };
    end 
    if(N1355) begin
      { data_buf_r[506:492] } <= { data_mem_data_i[506:492] };
    end 
    if(N1360) begin
      { data_buf_r[491:490] } <= { data_mem_data_i[491:490] };
    end 
    if(N1367) begin
      { data_buf_r[489:489] } <= { data_mem_data_i[489:489] };
    end 
    if(N1373) begin
      { data_buf_r[488:481] } <= { data_mem_data_i[488:481] };
    end 
    if(N1381) begin
      { data_buf_r[480:473] } <= { data_mem_data_i[480:473] };
    end 
    if(N1387) begin
      { data_buf_r[412:393] } <= { data_mem_data_i[412:393] };
    end 
    if(N1393) begin
      { data_buf_r[392:391] } <= { data_mem_data_i[392:391] };
    end 
    if(N1400) begin
      { data_buf_r[390:390] } <= { data_mem_data_i[390:390] };
    end 
    if(N1406) begin
      { data_buf_r[389:382] } <= { data_mem_data_i[389:382] };
    end 
    if(N1414) begin
      { data_buf_r[381:374] } <= { data_mem_data_i[381:374] };
    end 
    if(N1419) begin
      { data_buf_r[373:314] } <= { data_mem_data_i[373:314] };
    end 
    if(N1425) begin
      { data_buf_r[313:294] } <= { data_mem_data_i[313:294] };
    end 
    if(N1431) begin
      { data_buf_r[293:292] } <= { data_mem_data_i[293:292] };
    end 
    if(N1438) begin
      { data_buf_r[291:291] } <= { data_mem_data_i[291:291] };
    end 
    if(N1444) begin
      { data_buf_r[290:283] } <= { data_mem_data_i[290:283] };
    end 
    if(N1452) begin
      { data_buf_r[282:275] } <= { data_mem_data_i[282:275] };
    end 
    if(N1457) begin
      { data_buf_r[274:215] } <= { data_mem_data_i[274:215] };
    end 
    if(N1463) begin
      { data_buf_r[214:195] } <= { data_mem_data_i[214:195] };
    end 
    if(N1469) begin
      { data_buf_r[194:193] } <= { data_mem_data_i[194:193] };
    end 
    if(N1476) begin
      { data_buf_r[192:192] } <= { data_mem_data_i[192:192] };
    end 
    if(N1482) begin
      { data_buf_r[191:184] } <= { data_mem_data_i[191:184] };
    end 
    if(N1490) begin
      { data_buf_r[183:176] } <= { data_mem_data_i[183:176] };
    end 
    if(N1495) begin
      { data_buf_r[175:116] } <= { data_mem_data_i[175:116] };
    end 
    if(N1501) begin
      { data_buf_r[115:96] } <= { data_mem_data_i[115:96] };
    end 
    if(N1507) begin
      { data_buf_r[95:94] } <= { data_mem_data_i[95:94] };
    end 
    if(N1514) begin
      { data_buf_r[93:93] } <= { data_mem_data_i[93:93] };
    end 
    if(N1520) begin
      { data_buf_r[92:85] } <= { data_mem_data_i[92:85] };
    end 
    if(N1528) begin
      { data_buf_r[84:77] } <= { data_mem_data_i[84:77] };
    end 
    if(N1533) begin
      { data_buf_r[76:17], data_buf_r[4:4] } <= { data_mem_data_i[76:17], data_mem_data_i[4:4] };
    end 
    if(N1539) begin
      { data_buf_r[16:5] } <= { data_mem_data_i[16:5] };
    end 
    if(N1545) begin
      { data_buf_r[3:3] } <= { data_mem_data_i[3:3] };
    end 
    if(N1551) begin
      { data_buf_r[2:2] } <= { data_mem_data_i[2:2] };
    end 
    if(N1557) begin
      { data_buf_r[1:1] } <= { data_mem_data_i[1:1] };
    end 
    if(N1569) begin
      { state_r[2:0] } <= { N1247, N1246, N1245 };
    end 
    if(N1580) begin
      { sync_ack_count_r[0:0] } <= { N1248 };
    end 
    if(N1585) begin
      tr_data_buffered_r <= N1249;
    end 
    if(N1590) begin
      wb_data_buffered_r <= N1250;
      wb_data_read_r <= N1251;
      wb_dirty_cleared_r <= N1252;
    end 
    if(N1603) begin
      invalidated_tag_r <= N1253;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p540_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [539:0] w_data_i;
  input [0:0] r_addr_i;
  output [539:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [539:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  reg [1079:0] mem;
  assign r_data_o[539] = (N3)? mem[539] : 
                         (N0)? mem[1079] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[538] = (N3)? mem[538] : 
                         (N0)? mem[1078] : 1'b0;
  assign r_data_o[537] = (N3)? mem[537] : 
                         (N0)? mem[1077] : 1'b0;
  assign r_data_o[536] = (N3)? mem[536] : 
                         (N0)? mem[1076] : 1'b0;
  assign r_data_o[535] = (N3)? mem[535] : 
                         (N0)? mem[1075] : 1'b0;
  assign r_data_o[534] = (N3)? mem[534] : 
                         (N0)? mem[1074] : 1'b0;
  assign r_data_o[533] = (N3)? mem[533] : 
                         (N0)? mem[1073] : 1'b0;
  assign r_data_o[532] = (N3)? mem[532] : 
                         (N0)? mem[1072] : 1'b0;
  assign r_data_o[531] = (N3)? mem[531] : 
                         (N0)? mem[1071] : 1'b0;
  assign r_data_o[530] = (N3)? mem[530] : 
                         (N0)? mem[1070] : 1'b0;
  assign r_data_o[529] = (N3)? mem[529] : 
                         (N0)? mem[1069] : 1'b0;
  assign r_data_o[528] = (N3)? mem[528] : 
                         (N0)? mem[1068] : 1'b0;
  assign r_data_o[527] = (N3)? mem[527] : 
                         (N0)? mem[1067] : 1'b0;
  assign r_data_o[526] = (N3)? mem[526] : 
                         (N0)? mem[1066] : 1'b0;
  assign r_data_o[525] = (N3)? mem[525] : 
                         (N0)? mem[1065] : 1'b0;
  assign r_data_o[524] = (N3)? mem[524] : 
                         (N0)? mem[1064] : 1'b0;
  assign r_data_o[523] = (N3)? mem[523] : 
                         (N0)? mem[1063] : 1'b0;
  assign r_data_o[522] = (N3)? mem[522] : 
                         (N0)? mem[1062] : 1'b0;
  assign r_data_o[521] = (N3)? mem[521] : 
                         (N0)? mem[1061] : 1'b0;
  assign r_data_o[520] = (N3)? mem[520] : 
                         (N0)? mem[1060] : 1'b0;
  assign r_data_o[519] = (N3)? mem[519] : 
                         (N0)? mem[1059] : 1'b0;
  assign r_data_o[518] = (N3)? mem[518] : 
                         (N0)? mem[1058] : 1'b0;
  assign r_data_o[517] = (N3)? mem[517] : 
                         (N0)? mem[1057] : 1'b0;
  assign r_data_o[516] = (N3)? mem[516] : 
                         (N0)? mem[1056] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] : 
                         (N0)? mem[1055] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] : 
                         (N0)? mem[1054] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] : 
                         (N0)? mem[1053] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] : 
                         (N0)? mem[1052] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] : 
                         (N0)? mem[1051] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] : 
                         (N0)? mem[1050] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] : 
                         (N0)? mem[1049] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] : 
                         (N0)? mem[1048] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] : 
                         (N0)? mem[1047] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] : 
                         (N0)? mem[1046] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] : 
                         (N0)? mem[1045] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] : 
                         (N0)? mem[1044] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] : 
                         (N0)? mem[1043] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] : 
                         (N0)? mem[1042] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] : 
                         (N0)? mem[1041] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] : 
                         (N0)? mem[1040] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] : 
                         (N0)? mem[1039] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] : 
                         (N0)? mem[1038] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] : 
                         (N0)? mem[1037] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] : 
                         (N0)? mem[1036] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] : 
                         (N0)? mem[1035] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] : 
                         (N0)? mem[1034] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] : 
                         (N0)? mem[1033] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] : 
                         (N0)? mem[1032] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] : 
                         (N0)? mem[1031] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] : 
                         (N0)? mem[1030] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] : 
                         (N0)? mem[1029] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] : 
                         (N0)? mem[1028] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] : 
                         (N0)? mem[1027] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] : 
                         (N0)? mem[1026] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] : 
                         (N0)? mem[1025] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] : 
                         (N0)? mem[1024] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] : 
                         (N0)? mem[1023] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] : 
                         (N0)? mem[1022] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] : 
                         (N0)? mem[1021] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] : 
                         (N0)? mem[1020] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] : 
                         (N0)? mem[1019] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] : 
                         (N0)? mem[1018] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] : 
                         (N0)? mem[1017] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] : 
                         (N0)? mem[1016] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] : 
                         (N0)? mem[1015] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] : 
                         (N0)? mem[1014] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] : 
                         (N0)? mem[1013] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] : 
                         (N0)? mem[1012] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] : 
                         (N0)? mem[1011] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] : 
                         (N0)? mem[1010] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] : 
                         (N0)? mem[1009] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] : 
                         (N0)? mem[1008] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] : 
                         (N0)? mem[1007] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] : 
                         (N0)? mem[1006] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] : 
                         (N0)? mem[1005] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] : 
                         (N0)? mem[1004] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] : 
                         (N0)? mem[1003] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] : 
                         (N0)? mem[1002] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] : 
                         (N0)? mem[1001] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] : 
                         (N0)? mem[1000] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] : 
                         (N0)? mem[999] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] : 
                         (N0)? mem[998] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] : 
                         (N0)? mem[997] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] : 
                         (N0)? mem[996] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] : 
                         (N0)? mem[995] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] : 
                         (N0)? mem[994] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] : 
                         (N0)? mem[993] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] : 
                         (N0)? mem[992] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] : 
                         (N0)? mem[991] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] : 
                         (N0)? mem[990] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] : 
                         (N0)? mem[989] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] : 
                         (N0)? mem[988] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] : 
                         (N0)? mem[987] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] : 
                         (N0)? mem[986] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] : 
                         (N0)? mem[985] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] : 
                         (N0)? mem[984] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] : 
                         (N0)? mem[983] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] : 
                         (N0)? mem[982] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] : 
                         (N0)? mem[981] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] : 
                         (N0)? mem[980] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] : 
                         (N0)? mem[979] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] : 
                         (N0)? mem[978] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] : 
                         (N0)? mem[977] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] : 
                         (N0)? mem[976] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] : 
                         (N0)? mem[975] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] : 
                         (N0)? mem[974] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] : 
                         (N0)? mem[973] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] : 
                         (N0)? mem[972] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] : 
                         (N0)? mem[971] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] : 
                         (N0)? mem[970] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] : 
                         (N0)? mem[969] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] : 
                         (N0)? mem[968] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] : 
                         (N0)? mem[967] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] : 
                         (N0)? mem[966] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] : 
                         (N0)? mem[965] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] : 
                         (N0)? mem[964] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] : 
                         (N0)? mem[963] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] : 
                         (N0)? mem[962] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] : 
                         (N0)? mem[961] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] : 
                         (N0)? mem[960] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] : 
                         (N0)? mem[959] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] : 
                         (N0)? mem[958] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] : 
                         (N0)? mem[957] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] : 
                         (N0)? mem[956] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] : 
                         (N0)? mem[955] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] : 
                         (N0)? mem[954] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] : 
                         (N0)? mem[953] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] : 
                         (N0)? mem[952] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] : 
                         (N0)? mem[951] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] : 
                         (N0)? mem[950] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] : 
                         (N0)? mem[949] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] : 
                         (N0)? mem[948] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] : 
                         (N0)? mem[947] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] : 
                         (N0)? mem[946] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] : 
                         (N0)? mem[945] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] : 
                         (N0)? mem[944] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] : 
                         (N0)? mem[943] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] : 
                         (N0)? mem[942] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] : 
                         (N0)? mem[941] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] : 
                         (N0)? mem[940] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] : 
                         (N0)? mem[939] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] : 
                         (N0)? mem[938] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] : 
                         (N0)? mem[937] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] : 
                         (N0)? mem[936] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] : 
                         (N0)? mem[935] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] : 
                         (N0)? mem[934] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] : 
                         (N0)? mem[933] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] : 
                         (N0)? mem[932] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] : 
                         (N0)? mem[931] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] : 
                         (N0)? mem[930] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] : 
                         (N0)? mem[929] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] : 
                         (N0)? mem[928] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] : 
                         (N0)? mem[927] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] : 
                         (N0)? mem[926] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] : 
                         (N0)? mem[925] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] : 
                         (N0)? mem[924] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] : 
                         (N0)? mem[923] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] : 
                         (N0)? mem[922] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] : 
                         (N0)? mem[921] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] : 
                         (N0)? mem[920] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] : 
                         (N0)? mem[919] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] : 
                         (N0)? mem[918] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] : 
                         (N0)? mem[917] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] : 
                         (N0)? mem[916] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] : 
                         (N0)? mem[915] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] : 
                         (N0)? mem[914] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] : 
                         (N0)? mem[913] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] : 
                         (N0)? mem[912] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] : 
                         (N0)? mem[911] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] : 
                         (N0)? mem[910] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] : 
                         (N0)? mem[909] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] : 
                         (N0)? mem[908] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] : 
                         (N0)? mem[907] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] : 
                         (N0)? mem[906] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] : 
                         (N0)? mem[905] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] : 
                         (N0)? mem[904] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] : 
                         (N0)? mem[903] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] : 
                         (N0)? mem[902] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] : 
                         (N0)? mem[901] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] : 
                         (N0)? mem[900] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] : 
                         (N0)? mem[899] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] : 
                         (N0)? mem[898] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] : 
                         (N0)? mem[897] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] : 
                         (N0)? mem[896] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] : 
                         (N0)? mem[895] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] : 
                         (N0)? mem[894] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] : 
                         (N0)? mem[893] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] : 
                         (N0)? mem[892] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] : 
                         (N0)? mem[891] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] : 
                         (N0)? mem[890] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] : 
                         (N0)? mem[889] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] : 
                         (N0)? mem[888] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] : 
                         (N0)? mem[887] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] : 
                         (N0)? mem[886] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] : 
                         (N0)? mem[885] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] : 
                         (N0)? mem[884] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] : 
                         (N0)? mem[883] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] : 
                         (N0)? mem[882] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] : 
                         (N0)? mem[881] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] : 
                         (N0)? mem[880] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] : 
                         (N0)? mem[879] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] : 
                         (N0)? mem[878] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] : 
                         (N0)? mem[877] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] : 
                         (N0)? mem[876] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] : 
                         (N0)? mem[875] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] : 
                         (N0)? mem[874] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] : 
                         (N0)? mem[873] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] : 
                         (N0)? mem[872] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] : 
                         (N0)? mem[871] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] : 
                         (N0)? mem[870] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] : 
                         (N0)? mem[869] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] : 
                         (N0)? mem[868] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] : 
                         (N0)? mem[867] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] : 
                         (N0)? mem[866] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] : 
                         (N0)? mem[865] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] : 
                         (N0)? mem[864] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] : 
                         (N0)? mem[863] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] : 
                         (N0)? mem[862] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] : 
                         (N0)? mem[861] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] : 
                         (N0)? mem[860] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] : 
                         (N0)? mem[859] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] : 
                         (N0)? mem[858] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] : 
                         (N0)? mem[857] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] : 
                         (N0)? mem[856] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] : 
                         (N0)? mem[855] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] : 
                         (N0)? mem[854] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] : 
                         (N0)? mem[853] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] : 
                         (N0)? mem[852] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] : 
                         (N0)? mem[851] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] : 
                         (N0)? mem[850] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] : 
                         (N0)? mem[849] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] : 
                         (N0)? mem[848] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] : 
                         (N0)? mem[847] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] : 
                         (N0)? mem[846] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] : 
                         (N0)? mem[845] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] : 
                         (N0)? mem[844] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] : 
                         (N0)? mem[843] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] : 
                         (N0)? mem[842] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] : 
                         (N0)? mem[841] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] : 
                         (N0)? mem[840] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] : 
                         (N0)? mem[839] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] : 
                         (N0)? mem[838] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] : 
                         (N0)? mem[837] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] : 
                         (N0)? mem[836] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] : 
                         (N0)? mem[835] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] : 
                         (N0)? mem[834] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] : 
                         (N0)? mem[833] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] : 
                         (N0)? mem[832] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] : 
                         (N0)? mem[831] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] : 
                         (N0)? mem[830] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] : 
                         (N0)? mem[829] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] : 
                         (N0)? mem[828] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] : 
                         (N0)? mem[827] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] : 
                         (N0)? mem[826] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] : 
                         (N0)? mem[825] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] : 
                         (N0)? mem[824] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] : 
                         (N0)? mem[823] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] : 
                         (N0)? mem[822] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] : 
                         (N0)? mem[821] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] : 
                         (N0)? mem[820] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] : 
                         (N0)? mem[819] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] : 
                         (N0)? mem[818] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] : 
                         (N0)? mem[817] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] : 
                         (N0)? mem[816] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] : 
                         (N0)? mem[815] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] : 
                         (N0)? mem[814] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] : 
                         (N0)? mem[813] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] : 
                         (N0)? mem[812] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] : 
                         (N0)? mem[811] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] : 
                         (N0)? mem[810] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] : 
                         (N0)? mem[809] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] : 
                         (N0)? mem[808] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] : 
                         (N0)? mem[807] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] : 
                         (N0)? mem[806] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] : 
                         (N0)? mem[805] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] : 
                         (N0)? mem[804] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] : 
                         (N0)? mem[803] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] : 
                         (N0)? mem[802] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] : 
                         (N0)? mem[801] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] : 
                         (N0)? mem[800] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] : 
                         (N0)? mem[799] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] : 
                         (N0)? mem[798] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] : 
                         (N0)? mem[797] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] : 
                         (N0)? mem[796] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] : 
                         (N0)? mem[795] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] : 
                         (N0)? mem[794] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] : 
                         (N0)? mem[793] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] : 
                         (N0)? mem[792] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] : 
                         (N0)? mem[791] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] : 
                         (N0)? mem[790] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] : 
                         (N0)? mem[789] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] : 
                         (N0)? mem[788] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] : 
                         (N0)? mem[787] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] : 
                         (N0)? mem[786] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] : 
                         (N0)? mem[785] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] : 
                         (N0)? mem[784] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] : 
                         (N0)? mem[783] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] : 
                         (N0)? mem[782] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] : 
                         (N0)? mem[781] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] : 
                         (N0)? mem[780] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] : 
                         (N0)? mem[779] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] : 
                         (N0)? mem[778] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] : 
                         (N0)? mem[777] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] : 
                         (N0)? mem[776] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] : 
                         (N0)? mem[775] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] : 
                         (N0)? mem[774] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] : 
                         (N0)? mem[773] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] : 
                         (N0)? mem[772] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] : 
                         (N0)? mem[771] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] : 
                         (N0)? mem[770] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] : 
                         (N0)? mem[769] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] : 
                         (N0)? mem[768] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] : 
                         (N0)? mem[767] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] : 
                         (N0)? mem[766] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] : 
                         (N0)? mem[765] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] : 
                         (N0)? mem[764] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] : 
                         (N0)? mem[763] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] : 
                         (N0)? mem[762] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] : 
                         (N0)? mem[761] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] : 
                         (N0)? mem[760] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] : 
                         (N0)? mem[759] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] : 
                         (N0)? mem[758] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] : 
                         (N0)? mem[757] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] : 
                         (N0)? mem[756] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] : 
                         (N0)? mem[755] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] : 
                         (N0)? mem[754] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] : 
                         (N0)? mem[753] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] : 
                         (N0)? mem[752] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] : 
                         (N0)? mem[751] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] : 
                         (N0)? mem[750] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] : 
                         (N0)? mem[749] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] : 
                         (N0)? mem[748] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] : 
                         (N0)? mem[747] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] : 
                         (N0)? mem[746] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] : 
                         (N0)? mem[745] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] : 
                         (N0)? mem[744] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] : 
                         (N0)? mem[743] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] : 
                         (N0)? mem[742] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] : 
                         (N0)? mem[741] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] : 
                         (N0)? mem[740] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] : 
                         (N0)? mem[739] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] : 
                         (N0)? mem[738] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] : 
                         (N0)? mem[737] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] : 
                         (N0)? mem[736] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] : 
                         (N0)? mem[735] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] : 
                         (N0)? mem[734] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] : 
                         (N0)? mem[733] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] : 
                         (N0)? mem[732] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] : 
                         (N0)? mem[731] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] : 
                         (N0)? mem[730] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] : 
                         (N0)? mem[729] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] : 
                         (N0)? mem[728] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] : 
                         (N0)? mem[727] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] : 
                         (N0)? mem[726] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] : 
                         (N0)? mem[725] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] : 
                         (N0)? mem[724] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] : 
                         (N0)? mem[723] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] : 
                         (N0)? mem[722] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] : 
                         (N0)? mem[721] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] : 
                         (N0)? mem[720] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] : 
                         (N0)? mem[719] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] : 
                         (N0)? mem[718] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] : 
                         (N0)? mem[717] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] : 
                         (N0)? mem[716] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] : 
                         (N0)? mem[715] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] : 
                         (N0)? mem[714] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] : 
                         (N0)? mem[713] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] : 
                         (N0)? mem[712] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] : 
                         (N0)? mem[711] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] : 
                         (N0)? mem[710] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] : 
                         (N0)? mem[709] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] : 
                         (N0)? mem[708] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] : 
                         (N0)? mem[707] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] : 
                         (N0)? mem[706] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] : 
                         (N0)? mem[705] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] : 
                         (N0)? mem[704] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] : 
                         (N0)? mem[703] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] : 
                         (N0)? mem[702] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] : 
                         (N0)? mem[701] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] : 
                         (N0)? mem[700] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] : 
                         (N0)? mem[699] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] : 
                         (N0)? mem[698] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] : 
                         (N0)? mem[697] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] : 
                         (N0)? mem[696] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] : 
                         (N0)? mem[695] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] : 
                         (N0)? mem[694] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] : 
                         (N0)? mem[693] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] : 
                         (N0)? mem[692] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] : 
                         (N0)? mem[691] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] : 
                         (N0)? mem[690] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] : 
                         (N0)? mem[689] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] : 
                         (N0)? mem[688] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] : 
                         (N0)? mem[687] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] : 
                         (N0)? mem[686] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] : 
                         (N0)? mem[685] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] : 
                         (N0)? mem[684] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] : 
                         (N0)? mem[683] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] : 
                         (N0)? mem[682] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] : 
                         (N0)? mem[681] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] : 
                         (N0)? mem[680] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] : 
                         (N0)? mem[679] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] : 
                         (N0)? mem[678] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] : 
                         (N0)? mem[677] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] : 
                         (N0)? mem[676] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] : 
                         (N0)? mem[675] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] : 
                         (N0)? mem[674] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] : 
                         (N0)? mem[673] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] : 
                         (N0)? mem[672] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] : 
                         (N0)? mem[671] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] : 
                         (N0)? mem[670] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] : 
                         (N0)? mem[669] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] : 
                         (N0)? mem[668] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] : 
                         (N0)? mem[667] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] : 
                         (N0)? mem[666] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] : 
                         (N0)? mem[665] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] : 
                         (N0)? mem[664] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] : 
                         (N0)? mem[663] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] : 
                         (N0)? mem[662] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] : 
                         (N0)? mem[661] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] : 
                         (N0)? mem[660] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] : 
                         (N0)? mem[659] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] : 
                         (N0)? mem[658] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] : 
                         (N0)? mem[657] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] : 
                         (N0)? mem[656] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] : 
                         (N0)? mem[655] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] : 
                         (N0)? mem[654] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] : 
                         (N0)? mem[653] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] : 
                         (N0)? mem[652] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] : 
                         (N0)? mem[651] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] : 
                         (N0)? mem[650] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] : 
                         (N0)? mem[649] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] : 
                         (N0)? mem[648] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] : 
                         (N0)? mem[647] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] : 
                         (N0)? mem[646] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] : 
                         (N0)? mem[645] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] : 
                         (N0)? mem[644] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] : 
                         (N0)? mem[643] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] : 
                         (N0)? mem[642] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] : 
                         (N0)? mem[641] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] : 
                         (N0)? mem[640] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] : 
                        (N0)? mem[639] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] : 
                        (N0)? mem[638] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] : 
                        (N0)? mem[637] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] : 
                        (N0)? mem[636] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] : 
                        (N0)? mem[635] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] : 
                        (N0)? mem[634] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] : 
                        (N0)? mem[633] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] : 
                        (N0)? mem[632] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] : 
                        (N0)? mem[631] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] : 
                        (N0)? mem[630] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] : 
                        (N0)? mem[629] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] : 
                        (N0)? mem[628] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] : 
                        (N0)? mem[627] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] : 
                        (N0)? mem[626] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] : 
                        (N0)? mem[625] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] : 
                        (N0)? mem[624] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] : 
                        (N0)? mem[623] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] : 
                        (N0)? mem[622] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] : 
                        (N0)? mem[621] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] : 
                        (N0)? mem[620] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] : 
                        (N0)? mem[619] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] : 
                        (N0)? mem[618] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] : 
                        (N0)? mem[617] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] : 
                        (N0)? mem[616] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] : 
                        (N0)? mem[615] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] : 
                        (N0)? mem[614] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] : 
                        (N0)? mem[613] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] : 
                        (N0)? mem[612] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] : 
                        (N0)? mem[611] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] : 
                        (N0)? mem[610] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] : 
                        (N0)? mem[609] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] : 
                        (N0)? mem[608] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] : 
                        (N0)? mem[607] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] : 
                        (N0)? mem[606] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] : 
                        (N0)? mem[605] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] : 
                        (N0)? mem[604] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[603] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[602] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[601] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[600] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[599] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[598] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[597] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[596] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[595] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[594] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[593] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[592] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[591] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[590] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[589] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[588] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[587] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[586] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[585] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[584] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[583] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[582] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[581] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[580] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[579] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[578] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[577] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[576] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[575] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[574] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[573] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[572] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[571] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[570] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[569] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[568] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[567] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[566] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[565] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[564] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[563] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[562] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[561] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[560] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[559] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[558] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[557] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[556] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[555] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[554] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[553] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[552] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[551] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[550] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[549] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[548] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[547] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[546] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[545] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[544] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[543] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[542] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[541] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[540] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } : 
                                                                       (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N13) begin
      { mem[1079:981], mem[540:540] } <= { w_data_i[539:441], w_data_i[0:0] };
    end 
    if(N14) begin
      { mem[980:882], mem[541:541] } <= { w_data_i[440:342], w_data_i[1:1] };
    end 
    if(N15) begin
      { mem[881:783], mem[542:542] } <= { w_data_i[341:243], w_data_i[2:2] };
    end 
    if(N16) begin
      { mem[782:684], mem[543:543] } <= { w_data_i[242:144], w_data_i[3:3] };
    end 
    if(N17) begin
      { mem[683:585], mem[544:544] } <= { w_data_i[143:45], w_data_i[4:4] };
    end 
    if(N18) begin
      { mem[584:545] } <= { w_data_i[44:5] };
    end 
    if(N7) begin
      { mem[539:441], mem[0:0] } <= { w_data_i[539:441], w_data_i[0:0] };
    end 
    if(N8) begin
      { mem[440:342], mem[1:1] } <= { w_data_i[440:342], w_data_i[1:1] };
    end 
    if(N9) begin
      { mem[341:243], mem[2:2] } <= { w_data_i[341:243], w_data_i[2:2] };
    end 
    if(N10) begin
      { mem[242:144], mem[3:3] } <= { w_data_i[242:144], w_data_i[3:3] };
    end 
    if(N11) begin
      { mem[143:45], mem[4:4] } <= { w_data_i[143:45], w_data_i[4:4] };
    end 
    if(N12) begin
      { mem[44:5] } <= { w_data_i[44:5] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p540_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [539:0] w_data_i;
  input [0:0] r_addr_i;
  output [539:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [539:0] r_data_o;

  bsg_mem_1r1w_synth_width_p540_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p540
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [539:0] data_i;
  output [539:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [539:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p540_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bp_be_dcache_lce_data_cmd_num_cce_p1_num_lce_p2_data_width_p64_paddr_width_p22_lce_data_width_p512_ways_p8_sets_p64
(
  cce_data_received_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_yumi_o,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_pkt_yumi_i
);

  input [539:0] lce_data_cmd_i;
  output [521:0] data_mem_pkt_o;
  input lce_data_cmd_v_i;
  input data_mem_pkt_yumi_i;
  output cce_data_received_o;
  output lce_data_cmd_yumi_o;
  output data_mem_pkt_v_o;
  wire [521:0] data_mem_pkt_o;
  wire cce_data_received_o,lce_data_cmd_yumi_o,data_mem_pkt_v_o,data_mem_pkt_yumi_i,
  lce_data_cmd_v_i;
  assign data_mem_pkt_o[0] = 1'b1;
  assign cce_data_received_o = data_mem_pkt_yumi_i;
  assign lce_data_cmd_yumi_o = data_mem_pkt_yumi_i;
  assign data_mem_pkt_v_o = lce_data_cmd_v_i;
  assign data_mem_pkt_o[521] = lce_data_cmd_i[523];
  assign data_mem_pkt_o[520] = lce_data_cmd_i[522];
  assign data_mem_pkt_o[519] = lce_data_cmd_i[521];
  assign data_mem_pkt_o[518] = lce_data_cmd_i[520];
  assign data_mem_pkt_o[517] = lce_data_cmd_i[519];
  assign data_mem_pkt_o[516] = lce_data_cmd_i[518];
  assign data_mem_pkt_o[515] = lce_data_cmd_i[536];
  assign data_mem_pkt_o[514] = lce_data_cmd_i[535];
  assign data_mem_pkt_o[513] = lce_data_cmd_i[534];
  assign data_mem_pkt_o[512] = lce_data_cmd_i[511];
  assign data_mem_pkt_o[511] = lce_data_cmd_i[510];
  assign data_mem_pkt_o[510] = lce_data_cmd_i[509];
  assign data_mem_pkt_o[509] = lce_data_cmd_i[508];
  assign data_mem_pkt_o[508] = lce_data_cmd_i[507];
  assign data_mem_pkt_o[507] = lce_data_cmd_i[506];
  assign data_mem_pkt_o[506] = lce_data_cmd_i[505];
  assign data_mem_pkt_o[505] = lce_data_cmd_i[504];
  assign data_mem_pkt_o[504] = lce_data_cmd_i[503];
  assign data_mem_pkt_o[503] = lce_data_cmd_i[502];
  assign data_mem_pkt_o[502] = lce_data_cmd_i[501];
  assign data_mem_pkt_o[501] = lce_data_cmd_i[500];
  assign data_mem_pkt_o[500] = lce_data_cmd_i[499];
  assign data_mem_pkt_o[499] = lce_data_cmd_i[498];
  assign data_mem_pkt_o[498] = lce_data_cmd_i[497];
  assign data_mem_pkt_o[497] = lce_data_cmd_i[496];
  assign data_mem_pkt_o[496] = lce_data_cmd_i[495];
  assign data_mem_pkt_o[495] = lce_data_cmd_i[494];
  assign data_mem_pkt_o[494] = lce_data_cmd_i[493];
  assign data_mem_pkt_o[493] = lce_data_cmd_i[492];
  assign data_mem_pkt_o[492] = lce_data_cmd_i[491];
  assign data_mem_pkt_o[491] = lce_data_cmd_i[490];
  assign data_mem_pkt_o[490] = lce_data_cmd_i[489];
  assign data_mem_pkt_o[489] = lce_data_cmd_i[488];
  assign data_mem_pkt_o[488] = lce_data_cmd_i[487];
  assign data_mem_pkt_o[487] = lce_data_cmd_i[486];
  assign data_mem_pkt_o[486] = lce_data_cmd_i[485];
  assign data_mem_pkt_o[485] = lce_data_cmd_i[484];
  assign data_mem_pkt_o[484] = lce_data_cmd_i[483];
  assign data_mem_pkt_o[483] = lce_data_cmd_i[482];
  assign data_mem_pkt_o[482] = lce_data_cmd_i[481];
  assign data_mem_pkt_o[481] = lce_data_cmd_i[480];
  assign data_mem_pkt_o[480] = lce_data_cmd_i[479];
  assign data_mem_pkt_o[479] = lce_data_cmd_i[478];
  assign data_mem_pkt_o[478] = lce_data_cmd_i[477];
  assign data_mem_pkt_o[477] = lce_data_cmd_i[476];
  assign data_mem_pkt_o[476] = lce_data_cmd_i[475];
  assign data_mem_pkt_o[475] = lce_data_cmd_i[474];
  assign data_mem_pkt_o[474] = lce_data_cmd_i[473];
  assign data_mem_pkt_o[473] = lce_data_cmd_i[472];
  assign data_mem_pkt_o[472] = lce_data_cmd_i[471];
  assign data_mem_pkt_o[471] = lce_data_cmd_i[470];
  assign data_mem_pkt_o[470] = lce_data_cmd_i[469];
  assign data_mem_pkt_o[469] = lce_data_cmd_i[468];
  assign data_mem_pkt_o[468] = lce_data_cmd_i[467];
  assign data_mem_pkt_o[467] = lce_data_cmd_i[466];
  assign data_mem_pkt_o[466] = lce_data_cmd_i[465];
  assign data_mem_pkt_o[465] = lce_data_cmd_i[464];
  assign data_mem_pkt_o[464] = lce_data_cmd_i[463];
  assign data_mem_pkt_o[463] = lce_data_cmd_i[462];
  assign data_mem_pkt_o[462] = lce_data_cmd_i[461];
  assign data_mem_pkt_o[461] = lce_data_cmd_i[460];
  assign data_mem_pkt_o[460] = lce_data_cmd_i[459];
  assign data_mem_pkt_o[459] = lce_data_cmd_i[458];
  assign data_mem_pkt_o[458] = lce_data_cmd_i[457];
  assign data_mem_pkt_o[457] = lce_data_cmd_i[456];
  assign data_mem_pkt_o[456] = lce_data_cmd_i[455];
  assign data_mem_pkt_o[455] = lce_data_cmd_i[454];
  assign data_mem_pkt_o[454] = lce_data_cmd_i[453];
  assign data_mem_pkt_o[453] = lce_data_cmd_i[452];
  assign data_mem_pkt_o[452] = lce_data_cmd_i[451];
  assign data_mem_pkt_o[451] = lce_data_cmd_i[450];
  assign data_mem_pkt_o[450] = lce_data_cmd_i[449];
  assign data_mem_pkt_o[449] = lce_data_cmd_i[448];
  assign data_mem_pkt_o[448] = lce_data_cmd_i[447];
  assign data_mem_pkt_o[447] = lce_data_cmd_i[446];
  assign data_mem_pkt_o[446] = lce_data_cmd_i[445];
  assign data_mem_pkt_o[445] = lce_data_cmd_i[444];
  assign data_mem_pkt_o[444] = lce_data_cmd_i[443];
  assign data_mem_pkt_o[443] = lce_data_cmd_i[442];
  assign data_mem_pkt_o[442] = lce_data_cmd_i[441];
  assign data_mem_pkt_o[441] = lce_data_cmd_i[440];
  assign data_mem_pkt_o[440] = lce_data_cmd_i[439];
  assign data_mem_pkt_o[439] = lce_data_cmd_i[438];
  assign data_mem_pkt_o[438] = lce_data_cmd_i[437];
  assign data_mem_pkt_o[437] = lce_data_cmd_i[436];
  assign data_mem_pkt_o[436] = lce_data_cmd_i[435];
  assign data_mem_pkt_o[435] = lce_data_cmd_i[434];
  assign data_mem_pkt_o[434] = lce_data_cmd_i[433];
  assign data_mem_pkt_o[433] = lce_data_cmd_i[432];
  assign data_mem_pkt_o[432] = lce_data_cmd_i[431];
  assign data_mem_pkt_o[431] = lce_data_cmd_i[430];
  assign data_mem_pkt_o[430] = lce_data_cmd_i[429];
  assign data_mem_pkt_o[429] = lce_data_cmd_i[428];
  assign data_mem_pkt_o[428] = lce_data_cmd_i[427];
  assign data_mem_pkt_o[427] = lce_data_cmd_i[426];
  assign data_mem_pkt_o[426] = lce_data_cmd_i[425];
  assign data_mem_pkt_o[425] = lce_data_cmd_i[424];
  assign data_mem_pkt_o[424] = lce_data_cmd_i[423];
  assign data_mem_pkt_o[423] = lce_data_cmd_i[422];
  assign data_mem_pkt_o[422] = lce_data_cmd_i[421];
  assign data_mem_pkt_o[421] = lce_data_cmd_i[420];
  assign data_mem_pkt_o[420] = lce_data_cmd_i[419];
  assign data_mem_pkt_o[419] = lce_data_cmd_i[418];
  assign data_mem_pkt_o[418] = lce_data_cmd_i[417];
  assign data_mem_pkt_o[417] = lce_data_cmd_i[416];
  assign data_mem_pkt_o[416] = lce_data_cmd_i[415];
  assign data_mem_pkt_o[415] = lce_data_cmd_i[414];
  assign data_mem_pkt_o[414] = lce_data_cmd_i[413];
  assign data_mem_pkt_o[413] = lce_data_cmd_i[412];
  assign data_mem_pkt_o[412] = lce_data_cmd_i[411];
  assign data_mem_pkt_o[411] = lce_data_cmd_i[410];
  assign data_mem_pkt_o[410] = lce_data_cmd_i[409];
  assign data_mem_pkt_o[409] = lce_data_cmd_i[408];
  assign data_mem_pkt_o[408] = lce_data_cmd_i[407];
  assign data_mem_pkt_o[407] = lce_data_cmd_i[406];
  assign data_mem_pkt_o[406] = lce_data_cmd_i[405];
  assign data_mem_pkt_o[405] = lce_data_cmd_i[404];
  assign data_mem_pkt_o[404] = lce_data_cmd_i[403];
  assign data_mem_pkt_o[403] = lce_data_cmd_i[402];
  assign data_mem_pkt_o[402] = lce_data_cmd_i[401];
  assign data_mem_pkt_o[401] = lce_data_cmd_i[400];
  assign data_mem_pkt_o[400] = lce_data_cmd_i[399];
  assign data_mem_pkt_o[399] = lce_data_cmd_i[398];
  assign data_mem_pkt_o[398] = lce_data_cmd_i[397];
  assign data_mem_pkt_o[397] = lce_data_cmd_i[396];
  assign data_mem_pkt_o[396] = lce_data_cmd_i[395];
  assign data_mem_pkt_o[395] = lce_data_cmd_i[394];
  assign data_mem_pkt_o[394] = lce_data_cmd_i[393];
  assign data_mem_pkt_o[393] = lce_data_cmd_i[392];
  assign data_mem_pkt_o[392] = lce_data_cmd_i[391];
  assign data_mem_pkt_o[391] = lce_data_cmd_i[390];
  assign data_mem_pkt_o[390] = lce_data_cmd_i[389];
  assign data_mem_pkt_o[389] = lce_data_cmd_i[388];
  assign data_mem_pkt_o[388] = lce_data_cmd_i[387];
  assign data_mem_pkt_o[387] = lce_data_cmd_i[386];
  assign data_mem_pkt_o[386] = lce_data_cmd_i[385];
  assign data_mem_pkt_o[385] = lce_data_cmd_i[384];
  assign data_mem_pkt_o[384] = lce_data_cmd_i[383];
  assign data_mem_pkt_o[383] = lce_data_cmd_i[382];
  assign data_mem_pkt_o[382] = lce_data_cmd_i[381];
  assign data_mem_pkt_o[381] = lce_data_cmd_i[380];
  assign data_mem_pkt_o[380] = lce_data_cmd_i[379];
  assign data_mem_pkt_o[379] = lce_data_cmd_i[378];
  assign data_mem_pkt_o[378] = lce_data_cmd_i[377];
  assign data_mem_pkt_o[377] = lce_data_cmd_i[376];
  assign data_mem_pkt_o[376] = lce_data_cmd_i[375];
  assign data_mem_pkt_o[375] = lce_data_cmd_i[374];
  assign data_mem_pkt_o[374] = lce_data_cmd_i[373];
  assign data_mem_pkt_o[373] = lce_data_cmd_i[372];
  assign data_mem_pkt_o[372] = lce_data_cmd_i[371];
  assign data_mem_pkt_o[371] = lce_data_cmd_i[370];
  assign data_mem_pkt_o[370] = lce_data_cmd_i[369];
  assign data_mem_pkt_o[369] = lce_data_cmd_i[368];
  assign data_mem_pkt_o[368] = lce_data_cmd_i[367];
  assign data_mem_pkt_o[367] = lce_data_cmd_i[366];
  assign data_mem_pkt_o[366] = lce_data_cmd_i[365];
  assign data_mem_pkt_o[365] = lce_data_cmd_i[364];
  assign data_mem_pkt_o[364] = lce_data_cmd_i[363];
  assign data_mem_pkt_o[363] = lce_data_cmd_i[362];
  assign data_mem_pkt_o[362] = lce_data_cmd_i[361];
  assign data_mem_pkt_o[361] = lce_data_cmd_i[360];
  assign data_mem_pkt_o[360] = lce_data_cmd_i[359];
  assign data_mem_pkt_o[359] = lce_data_cmd_i[358];
  assign data_mem_pkt_o[358] = lce_data_cmd_i[357];
  assign data_mem_pkt_o[357] = lce_data_cmd_i[356];
  assign data_mem_pkt_o[356] = lce_data_cmd_i[355];
  assign data_mem_pkt_o[355] = lce_data_cmd_i[354];
  assign data_mem_pkt_o[354] = lce_data_cmd_i[353];
  assign data_mem_pkt_o[353] = lce_data_cmd_i[352];
  assign data_mem_pkt_o[352] = lce_data_cmd_i[351];
  assign data_mem_pkt_o[351] = lce_data_cmd_i[350];
  assign data_mem_pkt_o[350] = lce_data_cmd_i[349];
  assign data_mem_pkt_o[349] = lce_data_cmd_i[348];
  assign data_mem_pkt_o[348] = lce_data_cmd_i[347];
  assign data_mem_pkt_o[347] = lce_data_cmd_i[346];
  assign data_mem_pkt_o[346] = lce_data_cmd_i[345];
  assign data_mem_pkt_o[345] = lce_data_cmd_i[344];
  assign data_mem_pkt_o[344] = lce_data_cmd_i[343];
  assign data_mem_pkt_o[343] = lce_data_cmd_i[342];
  assign data_mem_pkt_o[342] = lce_data_cmd_i[341];
  assign data_mem_pkt_o[341] = lce_data_cmd_i[340];
  assign data_mem_pkt_o[340] = lce_data_cmd_i[339];
  assign data_mem_pkt_o[339] = lce_data_cmd_i[338];
  assign data_mem_pkt_o[338] = lce_data_cmd_i[337];
  assign data_mem_pkt_o[337] = lce_data_cmd_i[336];
  assign data_mem_pkt_o[336] = lce_data_cmd_i[335];
  assign data_mem_pkt_o[335] = lce_data_cmd_i[334];
  assign data_mem_pkt_o[334] = lce_data_cmd_i[333];
  assign data_mem_pkt_o[333] = lce_data_cmd_i[332];
  assign data_mem_pkt_o[332] = lce_data_cmd_i[331];
  assign data_mem_pkt_o[331] = lce_data_cmd_i[330];
  assign data_mem_pkt_o[330] = lce_data_cmd_i[329];
  assign data_mem_pkt_o[329] = lce_data_cmd_i[328];
  assign data_mem_pkt_o[328] = lce_data_cmd_i[327];
  assign data_mem_pkt_o[327] = lce_data_cmd_i[326];
  assign data_mem_pkt_o[326] = lce_data_cmd_i[325];
  assign data_mem_pkt_o[325] = lce_data_cmd_i[324];
  assign data_mem_pkt_o[324] = lce_data_cmd_i[323];
  assign data_mem_pkt_o[323] = lce_data_cmd_i[322];
  assign data_mem_pkt_o[322] = lce_data_cmd_i[321];
  assign data_mem_pkt_o[321] = lce_data_cmd_i[320];
  assign data_mem_pkt_o[320] = lce_data_cmd_i[319];
  assign data_mem_pkt_o[319] = lce_data_cmd_i[318];
  assign data_mem_pkt_o[318] = lce_data_cmd_i[317];
  assign data_mem_pkt_o[317] = lce_data_cmd_i[316];
  assign data_mem_pkt_o[316] = lce_data_cmd_i[315];
  assign data_mem_pkt_o[315] = lce_data_cmd_i[314];
  assign data_mem_pkt_o[314] = lce_data_cmd_i[313];
  assign data_mem_pkt_o[313] = lce_data_cmd_i[312];
  assign data_mem_pkt_o[312] = lce_data_cmd_i[311];
  assign data_mem_pkt_o[311] = lce_data_cmd_i[310];
  assign data_mem_pkt_o[310] = lce_data_cmd_i[309];
  assign data_mem_pkt_o[309] = lce_data_cmd_i[308];
  assign data_mem_pkt_o[308] = lce_data_cmd_i[307];
  assign data_mem_pkt_o[307] = lce_data_cmd_i[306];
  assign data_mem_pkt_o[306] = lce_data_cmd_i[305];
  assign data_mem_pkt_o[305] = lce_data_cmd_i[304];
  assign data_mem_pkt_o[304] = lce_data_cmd_i[303];
  assign data_mem_pkt_o[303] = lce_data_cmd_i[302];
  assign data_mem_pkt_o[302] = lce_data_cmd_i[301];
  assign data_mem_pkt_o[301] = lce_data_cmd_i[300];
  assign data_mem_pkt_o[300] = lce_data_cmd_i[299];
  assign data_mem_pkt_o[299] = lce_data_cmd_i[298];
  assign data_mem_pkt_o[298] = lce_data_cmd_i[297];
  assign data_mem_pkt_o[297] = lce_data_cmd_i[296];
  assign data_mem_pkt_o[296] = lce_data_cmd_i[295];
  assign data_mem_pkt_o[295] = lce_data_cmd_i[294];
  assign data_mem_pkt_o[294] = lce_data_cmd_i[293];
  assign data_mem_pkt_o[293] = lce_data_cmd_i[292];
  assign data_mem_pkt_o[292] = lce_data_cmd_i[291];
  assign data_mem_pkt_o[291] = lce_data_cmd_i[290];
  assign data_mem_pkt_o[290] = lce_data_cmd_i[289];
  assign data_mem_pkt_o[289] = lce_data_cmd_i[288];
  assign data_mem_pkt_o[288] = lce_data_cmd_i[287];
  assign data_mem_pkt_o[287] = lce_data_cmd_i[286];
  assign data_mem_pkt_o[286] = lce_data_cmd_i[285];
  assign data_mem_pkt_o[285] = lce_data_cmd_i[284];
  assign data_mem_pkt_o[284] = lce_data_cmd_i[283];
  assign data_mem_pkt_o[283] = lce_data_cmd_i[282];
  assign data_mem_pkt_o[282] = lce_data_cmd_i[281];
  assign data_mem_pkt_o[281] = lce_data_cmd_i[280];
  assign data_mem_pkt_o[280] = lce_data_cmd_i[279];
  assign data_mem_pkt_o[279] = lce_data_cmd_i[278];
  assign data_mem_pkt_o[278] = lce_data_cmd_i[277];
  assign data_mem_pkt_o[277] = lce_data_cmd_i[276];
  assign data_mem_pkt_o[276] = lce_data_cmd_i[275];
  assign data_mem_pkt_o[275] = lce_data_cmd_i[274];
  assign data_mem_pkt_o[274] = lce_data_cmd_i[273];
  assign data_mem_pkt_o[273] = lce_data_cmd_i[272];
  assign data_mem_pkt_o[272] = lce_data_cmd_i[271];
  assign data_mem_pkt_o[271] = lce_data_cmd_i[270];
  assign data_mem_pkt_o[270] = lce_data_cmd_i[269];
  assign data_mem_pkt_o[269] = lce_data_cmd_i[268];
  assign data_mem_pkt_o[268] = lce_data_cmd_i[267];
  assign data_mem_pkt_o[267] = lce_data_cmd_i[266];
  assign data_mem_pkt_o[266] = lce_data_cmd_i[265];
  assign data_mem_pkt_o[265] = lce_data_cmd_i[264];
  assign data_mem_pkt_o[264] = lce_data_cmd_i[263];
  assign data_mem_pkt_o[263] = lce_data_cmd_i[262];
  assign data_mem_pkt_o[262] = lce_data_cmd_i[261];
  assign data_mem_pkt_o[261] = lce_data_cmd_i[260];
  assign data_mem_pkt_o[260] = lce_data_cmd_i[259];
  assign data_mem_pkt_o[259] = lce_data_cmd_i[258];
  assign data_mem_pkt_o[258] = lce_data_cmd_i[257];
  assign data_mem_pkt_o[257] = lce_data_cmd_i[256];
  assign data_mem_pkt_o[256] = lce_data_cmd_i[255];
  assign data_mem_pkt_o[255] = lce_data_cmd_i[254];
  assign data_mem_pkt_o[254] = lce_data_cmd_i[253];
  assign data_mem_pkt_o[253] = lce_data_cmd_i[252];
  assign data_mem_pkt_o[252] = lce_data_cmd_i[251];
  assign data_mem_pkt_o[251] = lce_data_cmd_i[250];
  assign data_mem_pkt_o[250] = lce_data_cmd_i[249];
  assign data_mem_pkt_o[249] = lce_data_cmd_i[248];
  assign data_mem_pkt_o[248] = lce_data_cmd_i[247];
  assign data_mem_pkt_o[247] = lce_data_cmd_i[246];
  assign data_mem_pkt_o[246] = lce_data_cmd_i[245];
  assign data_mem_pkt_o[245] = lce_data_cmd_i[244];
  assign data_mem_pkt_o[244] = lce_data_cmd_i[243];
  assign data_mem_pkt_o[243] = lce_data_cmd_i[242];
  assign data_mem_pkt_o[242] = lce_data_cmd_i[241];
  assign data_mem_pkt_o[241] = lce_data_cmd_i[240];
  assign data_mem_pkt_o[240] = lce_data_cmd_i[239];
  assign data_mem_pkt_o[239] = lce_data_cmd_i[238];
  assign data_mem_pkt_o[238] = lce_data_cmd_i[237];
  assign data_mem_pkt_o[237] = lce_data_cmd_i[236];
  assign data_mem_pkt_o[236] = lce_data_cmd_i[235];
  assign data_mem_pkt_o[235] = lce_data_cmd_i[234];
  assign data_mem_pkt_o[234] = lce_data_cmd_i[233];
  assign data_mem_pkt_o[233] = lce_data_cmd_i[232];
  assign data_mem_pkt_o[232] = lce_data_cmd_i[231];
  assign data_mem_pkt_o[231] = lce_data_cmd_i[230];
  assign data_mem_pkt_o[230] = lce_data_cmd_i[229];
  assign data_mem_pkt_o[229] = lce_data_cmd_i[228];
  assign data_mem_pkt_o[228] = lce_data_cmd_i[227];
  assign data_mem_pkt_o[227] = lce_data_cmd_i[226];
  assign data_mem_pkt_o[226] = lce_data_cmd_i[225];
  assign data_mem_pkt_o[225] = lce_data_cmd_i[224];
  assign data_mem_pkt_o[224] = lce_data_cmd_i[223];
  assign data_mem_pkt_o[223] = lce_data_cmd_i[222];
  assign data_mem_pkt_o[222] = lce_data_cmd_i[221];
  assign data_mem_pkt_o[221] = lce_data_cmd_i[220];
  assign data_mem_pkt_o[220] = lce_data_cmd_i[219];
  assign data_mem_pkt_o[219] = lce_data_cmd_i[218];
  assign data_mem_pkt_o[218] = lce_data_cmd_i[217];
  assign data_mem_pkt_o[217] = lce_data_cmd_i[216];
  assign data_mem_pkt_o[216] = lce_data_cmd_i[215];
  assign data_mem_pkt_o[215] = lce_data_cmd_i[214];
  assign data_mem_pkt_o[214] = lce_data_cmd_i[213];
  assign data_mem_pkt_o[213] = lce_data_cmd_i[212];
  assign data_mem_pkt_o[212] = lce_data_cmd_i[211];
  assign data_mem_pkt_o[211] = lce_data_cmd_i[210];
  assign data_mem_pkt_o[210] = lce_data_cmd_i[209];
  assign data_mem_pkt_o[209] = lce_data_cmd_i[208];
  assign data_mem_pkt_o[208] = lce_data_cmd_i[207];
  assign data_mem_pkt_o[207] = lce_data_cmd_i[206];
  assign data_mem_pkt_o[206] = lce_data_cmd_i[205];
  assign data_mem_pkt_o[205] = lce_data_cmd_i[204];
  assign data_mem_pkt_o[204] = lce_data_cmd_i[203];
  assign data_mem_pkt_o[203] = lce_data_cmd_i[202];
  assign data_mem_pkt_o[202] = lce_data_cmd_i[201];
  assign data_mem_pkt_o[201] = lce_data_cmd_i[200];
  assign data_mem_pkt_o[200] = lce_data_cmd_i[199];
  assign data_mem_pkt_o[199] = lce_data_cmd_i[198];
  assign data_mem_pkt_o[198] = lce_data_cmd_i[197];
  assign data_mem_pkt_o[197] = lce_data_cmd_i[196];
  assign data_mem_pkt_o[196] = lce_data_cmd_i[195];
  assign data_mem_pkt_o[195] = lce_data_cmd_i[194];
  assign data_mem_pkt_o[194] = lce_data_cmd_i[193];
  assign data_mem_pkt_o[193] = lce_data_cmd_i[192];
  assign data_mem_pkt_o[192] = lce_data_cmd_i[191];
  assign data_mem_pkt_o[191] = lce_data_cmd_i[190];
  assign data_mem_pkt_o[190] = lce_data_cmd_i[189];
  assign data_mem_pkt_o[189] = lce_data_cmd_i[188];
  assign data_mem_pkt_o[188] = lce_data_cmd_i[187];
  assign data_mem_pkt_o[187] = lce_data_cmd_i[186];
  assign data_mem_pkt_o[186] = lce_data_cmd_i[185];
  assign data_mem_pkt_o[185] = lce_data_cmd_i[184];
  assign data_mem_pkt_o[184] = lce_data_cmd_i[183];
  assign data_mem_pkt_o[183] = lce_data_cmd_i[182];
  assign data_mem_pkt_o[182] = lce_data_cmd_i[181];
  assign data_mem_pkt_o[181] = lce_data_cmd_i[180];
  assign data_mem_pkt_o[180] = lce_data_cmd_i[179];
  assign data_mem_pkt_o[179] = lce_data_cmd_i[178];
  assign data_mem_pkt_o[178] = lce_data_cmd_i[177];
  assign data_mem_pkt_o[177] = lce_data_cmd_i[176];
  assign data_mem_pkt_o[176] = lce_data_cmd_i[175];
  assign data_mem_pkt_o[175] = lce_data_cmd_i[174];
  assign data_mem_pkt_o[174] = lce_data_cmd_i[173];
  assign data_mem_pkt_o[173] = lce_data_cmd_i[172];
  assign data_mem_pkt_o[172] = lce_data_cmd_i[171];
  assign data_mem_pkt_o[171] = lce_data_cmd_i[170];
  assign data_mem_pkt_o[170] = lce_data_cmd_i[169];
  assign data_mem_pkt_o[169] = lce_data_cmd_i[168];
  assign data_mem_pkt_o[168] = lce_data_cmd_i[167];
  assign data_mem_pkt_o[167] = lce_data_cmd_i[166];
  assign data_mem_pkt_o[166] = lce_data_cmd_i[165];
  assign data_mem_pkt_o[165] = lce_data_cmd_i[164];
  assign data_mem_pkt_o[164] = lce_data_cmd_i[163];
  assign data_mem_pkt_o[163] = lce_data_cmd_i[162];
  assign data_mem_pkt_o[162] = lce_data_cmd_i[161];
  assign data_mem_pkt_o[161] = lce_data_cmd_i[160];
  assign data_mem_pkt_o[160] = lce_data_cmd_i[159];
  assign data_mem_pkt_o[159] = lce_data_cmd_i[158];
  assign data_mem_pkt_o[158] = lce_data_cmd_i[157];
  assign data_mem_pkt_o[157] = lce_data_cmd_i[156];
  assign data_mem_pkt_o[156] = lce_data_cmd_i[155];
  assign data_mem_pkt_o[155] = lce_data_cmd_i[154];
  assign data_mem_pkt_o[154] = lce_data_cmd_i[153];
  assign data_mem_pkt_o[153] = lce_data_cmd_i[152];
  assign data_mem_pkt_o[152] = lce_data_cmd_i[151];
  assign data_mem_pkt_o[151] = lce_data_cmd_i[150];
  assign data_mem_pkt_o[150] = lce_data_cmd_i[149];
  assign data_mem_pkt_o[149] = lce_data_cmd_i[148];
  assign data_mem_pkt_o[148] = lce_data_cmd_i[147];
  assign data_mem_pkt_o[147] = lce_data_cmd_i[146];
  assign data_mem_pkt_o[146] = lce_data_cmd_i[145];
  assign data_mem_pkt_o[145] = lce_data_cmd_i[144];
  assign data_mem_pkt_o[144] = lce_data_cmd_i[143];
  assign data_mem_pkt_o[143] = lce_data_cmd_i[142];
  assign data_mem_pkt_o[142] = lce_data_cmd_i[141];
  assign data_mem_pkt_o[141] = lce_data_cmd_i[140];
  assign data_mem_pkt_o[140] = lce_data_cmd_i[139];
  assign data_mem_pkt_o[139] = lce_data_cmd_i[138];
  assign data_mem_pkt_o[138] = lce_data_cmd_i[137];
  assign data_mem_pkt_o[137] = lce_data_cmd_i[136];
  assign data_mem_pkt_o[136] = lce_data_cmd_i[135];
  assign data_mem_pkt_o[135] = lce_data_cmd_i[134];
  assign data_mem_pkt_o[134] = lce_data_cmd_i[133];
  assign data_mem_pkt_o[133] = lce_data_cmd_i[132];
  assign data_mem_pkt_o[132] = lce_data_cmd_i[131];
  assign data_mem_pkt_o[131] = lce_data_cmd_i[130];
  assign data_mem_pkt_o[130] = lce_data_cmd_i[129];
  assign data_mem_pkt_o[129] = lce_data_cmd_i[128];
  assign data_mem_pkt_o[128] = lce_data_cmd_i[127];
  assign data_mem_pkt_o[127] = lce_data_cmd_i[126];
  assign data_mem_pkt_o[126] = lce_data_cmd_i[125];
  assign data_mem_pkt_o[125] = lce_data_cmd_i[124];
  assign data_mem_pkt_o[124] = lce_data_cmd_i[123];
  assign data_mem_pkt_o[123] = lce_data_cmd_i[122];
  assign data_mem_pkt_o[122] = lce_data_cmd_i[121];
  assign data_mem_pkt_o[121] = lce_data_cmd_i[120];
  assign data_mem_pkt_o[120] = lce_data_cmd_i[119];
  assign data_mem_pkt_o[119] = lce_data_cmd_i[118];
  assign data_mem_pkt_o[118] = lce_data_cmd_i[117];
  assign data_mem_pkt_o[117] = lce_data_cmd_i[116];
  assign data_mem_pkt_o[116] = lce_data_cmd_i[115];
  assign data_mem_pkt_o[115] = lce_data_cmd_i[114];
  assign data_mem_pkt_o[114] = lce_data_cmd_i[113];
  assign data_mem_pkt_o[113] = lce_data_cmd_i[112];
  assign data_mem_pkt_o[112] = lce_data_cmd_i[111];
  assign data_mem_pkt_o[111] = lce_data_cmd_i[110];
  assign data_mem_pkt_o[110] = lce_data_cmd_i[109];
  assign data_mem_pkt_o[109] = lce_data_cmd_i[108];
  assign data_mem_pkt_o[108] = lce_data_cmd_i[107];
  assign data_mem_pkt_o[107] = lce_data_cmd_i[106];
  assign data_mem_pkt_o[106] = lce_data_cmd_i[105];
  assign data_mem_pkt_o[105] = lce_data_cmd_i[104];
  assign data_mem_pkt_o[104] = lce_data_cmd_i[103];
  assign data_mem_pkt_o[103] = lce_data_cmd_i[102];
  assign data_mem_pkt_o[102] = lce_data_cmd_i[101];
  assign data_mem_pkt_o[101] = lce_data_cmd_i[100];
  assign data_mem_pkt_o[100] = lce_data_cmd_i[99];
  assign data_mem_pkt_o[99] = lce_data_cmd_i[98];
  assign data_mem_pkt_o[98] = lce_data_cmd_i[97];
  assign data_mem_pkt_o[97] = lce_data_cmd_i[96];
  assign data_mem_pkt_o[96] = lce_data_cmd_i[95];
  assign data_mem_pkt_o[95] = lce_data_cmd_i[94];
  assign data_mem_pkt_o[94] = lce_data_cmd_i[93];
  assign data_mem_pkt_o[93] = lce_data_cmd_i[92];
  assign data_mem_pkt_o[92] = lce_data_cmd_i[91];
  assign data_mem_pkt_o[91] = lce_data_cmd_i[90];
  assign data_mem_pkt_o[90] = lce_data_cmd_i[89];
  assign data_mem_pkt_o[89] = lce_data_cmd_i[88];
  assign data_mem_pkt_o[88] = lce_data_cmd_i[87];
  assign data_mem_pkt_o[87] = lce_data_cmd_i[86];
  assign data_mem_pkt_o[86] = lce_data_cmd_i[85];
  assign data_mem_pkt_o[85] = lce_data_cmd_i[84];
  assign data_mem_pkt_o[84] = lce_data_cmd_i[83];
  assign data_mem_pkt_o[83] = lce_data_cmd_i[82];
  assign data_mem_pkt_o[82] = lce_data_cmd_i[81];
  assign data_mem_pkt_o[81] = lce_data_cmd_i[80];
  assign data_mem_pkt_o[80] = lce_data_cmd_i[79];
  assign data_mem_pkt_o[79] = lce_data_cmd_i[78];
  assign data_mem_pkt_o[78] = lce_data_cmd_i[77];
  assign data_mem_pkt_o[77] = lce_data_cmd_i[76];
  assign data_mem_pkt_o[76] = lce_data_cmd_i[75];
  assign data_mem_pkt_o[75] = lce_data_cmd_i[74];
  assign data_mem_pkt_o[74] = lce_data_cmd_i[73];
  assign data_mem_pkt_o[73] = lce_data_cmd_i[72];
  assign data_mem_pkt_o[72] = lce_data_cmd_i[71];
  assign data_mem_pkt_o[71] = lce_data_cmd_i[70];
  assign data_mem_pkt_o[70] = lce_data_cmd_i[69];
  assign data_mem_pkt_o[69] = lce_data_cmd_i[68];
  assign data_mem_pkt_o[68] = lce_data_cmd_i[67];
  assign data_mem_pkt_o[67] = lce_data_cmd_i[66];
  assign data_mem_pkt_o[66] = lce_data_cmd_i[65];
  assign data_mem_pkt_o[65] = lce_data_cmd_i[64];
  assign data_mem_pkt_o[64] = lce_data_cmd_i[63];
  assign data_mem_pkt_o[63] = lce_data_cmd_i[62];
  assign data_mem_pkt_o[62] = lce_data_cmd_i[61];
  assign data_mem_pkt_o[61] = lce_data_cmd_i[60];
  assign data_mem_pkt_o[60] = lce_data_cmd_i[59];
  assign data_mem_pkt_o[59] = lce_data_cmd_i[58];
  assign data_mem_pkt_o[58] = lce_data_cmd_i[57];
  assign data_mem_pkt_o[57] = lce_data_cmd_i[56];
  assign data_mem_pkt_o[56] = lce_data_cmd_i[55];
  assign data_mem_pkt_o[55] = lce_data_cmd_i[54];
  assign data_mem_pkt_o[54] = lce_data_cmd_i[53];
  assign data_mem_pkt_o[53] = lce_data_cmd_i[52];
  assign data_mem_pkt_o[52] = lce_data_cmd_i[51];
  assign data_mem_pkt_o[51] = lce_data_cmd_i[50];
  assign data_mem_pkt_o[50] = lce_data_cmd_i[49];
  assign data_mem_pkt_o[49] = lce_data_cmd_i[48];
  assign data_mem_pkt_o[48] = lce_data_cmd_i[47];
  assign data_mem_pkt_o[47] = lce_data_cmd_i[46];
  assign data_mem_pkt_o[46] = lce_data_cmd_i[45];
  assign data_mem_pkt_o[45] = lce_data_cmd_i[44];
  assign data_mem_pkt_o[44] = lce_data_cmd_i[43];
  assign data_mem_pkt_o[43] = lce_data_cmd_i[42];
  assign data_mem_pkt_o[42] = lce_data_cmd_i[41];
  assign data_mem_pkt_o[41] = lce_data_cmd_i[40];
  assign data_mem_pkt_o[40] = lce_data_cmd_i[39];
  assign data_mem_pkt_o[39] = lce_data_cmd_i[38];
  assign data_mem_pkt_o[38] = lce_data_cmd_i[37];
  assign data_mem_pkt_o[37] = lce_data_cmd_i[36];
  assign data_mem_pkt_o[36] = lce_data_cmd_i[35];
  assign data_mem_pkt_o[35] = lce_data_cmd_i[34];
  assign data_mem_pkt_o[34] = lce_data_cmd_i[33];
  assign data_mem_pkt_o[33] = lce_data_cmd_i[32];
  assign data_mem_pkt_o[32] = lce_data_cmd_i[31];
  assign data_mem_pkt_o[31] = lce_data_cmd_i[30];
  assign data_mem_pkt_o[30] = lce_data_cmd_i[29];
  assign data_mem_pkt_o[29] = lce_data_cmd_i[28];
  assign data_mem_pkt_o[28] = lce_data_cmd_i[27];
  assign data_mem_pkt_o[27] = lce_data_cmd_i[26];
  assign data_mem_pkt_o[26] = lce_data_cmd_i[25];
  assign data_mem_pkt_o[25] = lce_data_cmd_i[24];
  assign data_mem_pkt_o[24] = lce_data_cmd_i[23];
  assign data_mem_pkt_o[23] = lce_data_cmd_i[22];
  assign data_mem_pkt_o[22] = lce_data_cmd_i[21];
  assign data_mem_pkt_o[21] = lce_data_cmd_i[20];
  assign data_mem_pkt_o[20] = lce_data_cmd_i[19];
  assign data_mem_pkt_o[19] = lce_data_cmd_i[18];
  assign data_mem_pkt_o[18] = lce_data_cmd_i[17];
  assign data_mem_pkt_o[17] = lce_data_cmd_i[16];
  assign data_mem_pkt_o[16] = lce_data_cmd_i[15];
  assign data_mem_pkt_o[15] = lce_data_cmd_i[14];
  assign data_mem_pkt_o[14] = lce_data_cmd_i[13];
  assign data_mem_pkt_o[13] = lce_data_cmd_i[12];
  assign data_mem_pkt_o[12] = lce_data_cmd_i[11];
  assign data_mem_pkt_o[11] = lce_data_cmd_i[10];
  assign data_mem_pkt_o[10] = lce_data_cmd_i[9];
  assign data_mem_pkt_o[9] = lce_data_cmd_i[8];
  assign data_mem_pkt_o[8] = lce_data_cmd_i[7];
  assign data_mem_pkt_o[7] = lce_data_cmd_i[6];
  assign data_mem_pkt_o[6] = lce_data_cmd_i[5];
  assign data_mem_pkt_o[5] = lce_data_cmd_i[4];
  assign data_mem_pkt_o[4] = lce_data_cmd_i[3];
  assign data_mem_pkt_o[3] = lce_data_cmd_i[2];
  assign data_mem_pkt_o[2] = lce_data_cmd_i[1];
  assign data_mem_pkt_o[1] = lce_data_cmd_i[0];

endmodule



module bsg_mem_1r1w_synth_width_p539_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [538:0] w_data_i;
  input [0:0] r_addr_i;
  output [538:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [538:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  reg [1077:0] mem;
  assign r_data_o[538] = (N3)? mem[538] : 
                         (N0)? mem[1077] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[537] = (N3)? mem[537] : 
                         (N0)? mem[1076] : 1'b0;
  assign r_data_o[536] = (N3)? mem[536] : 
                         (N0)? mem[1075] : 1'b0;
  assign r_data_o[535] = (N3)? mem[535] : 
                         (N0)? mem[1074] : 1'b0;
  assign r_data_o[534] = (N3)? mem[534] : 
                         (N0)? mem[1073] : 1'b0;
  assign r_data_o[533] = (N3)? mem[533] : 
                         (N0)? mem[1072] : 1'b0;
  assign r_data_o[532] = (N3)? mem[532] : 
                         (N0)? mem[1071] : 1'b0;
  assign r_data_o[531] = (N3)? mem[531] : 
                         (N0)? mem[1070] : 1'b0;
  assign r_data_o[530] = (N3)? mem[530] : 
                         (N0)? mem[1069] : 1'b0;
  assign r_data_o[529] = (N3)? mem[529] : 
                         (N0)? mem[1068] : 1'b0;
  assign r_data_o[528] = (N3)? mem[528] : 
                         (N0)? mem[1067] : 1'b0;
  assign r_data_o[527] = (N3)? mem[527] : 
                         (N0)? mem[1066] : 1'b0;
  assign r_data_o[526] = (N3)? mem[526] : 
                         (N0)? mem[1065] : 1'b0;
  assign r_data_o[525] = (N3)? mem[525] : 
                         (N0)? mem[1064] : 1'b0;
  assign r_data_o[524] = (N3)? mem[524] : 
                         (N0)? mem[1063] : 1'b0;
  assign r_data_o[523] = (N3)? mem[523] : 
                         (N0)? mem[1062] : 1'b0;
  assign r_data_o[522] = (N3)? mem[522] : 
                         (N0)? mem[1061] : 1'b0;
  assign r_data_o[521] = (N3)? mem[521] : 
                         (N0)? mem[1060] : 1'b0;
  assign r_data_o[520] = (N3)? mem[520] : 
                         (N0)? mem[1059] : 1'b0;
  assign r_data_o[519] = (N3)? mem[519] : 
                         (N0)? mem[1058] : 1'b0;
  assign r_data_o[518] = (N3)? mem[518] : 
                         (N0)? mem[1057] : 1'b0;
  assign r_data_o[517] = (N3)? mem[517] : 
                         (N0)? mem[1056] : 1'b0;
  assign r_data_o[516] = (N3)? mem[516] : 
                         (N0)? mem[1055] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] : 
                         (N0)? mem[1054] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] : 
                         (N0)? mem[1053] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] : 
                         (N0)? mem[1052] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] : 
                         (N0)? mem[1051] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] : 
                         (N0)? mem[1050] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] : 
                         (N0)? mem[1049] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] : 
                         (N0)? mem[1048] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] : 
                         (N0)? mem[1047] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] : 
                         (N0)? mem[1046] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] : 
                         (N0)? mem[1045] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] : 
                         (N0)? mem[1044] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] : 
                         (N0)? mem[1043] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] : 
                         (N0)? mem[1042] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] : 
                         (N0)? mem[1041] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] : 
                         (N0)? mem[1040] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] : 
                         (N0)? mem[1039] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] : 
                         (N0)? mem[1038] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] : 
                         (N0)? mem[1037] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] : 
                         (N0)? mem[1036] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] : 
                         (N0)? mem[1035] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] : 
                         (N0)? mem[1034] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] : 
                         (N0)? mem[1033] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] : 
                         (N0)? mem[1032] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] : 
                         (N0)? mem[1031] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] : 
                         (N0)? mem[1030] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] : 
                         (N0)? mem[1029] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] : 
                         (N0)? mem[1028] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] : 
                         (N0)? mem[1027] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] : 
                         (N0)? mem[1026] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] : 
                         (N0)? mem[1025] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] : 
                         (N0)? mem[1024] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] : 
                         (N0)? mem[1023] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] : 
                         (N0)? mem[1022] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] : 
                         (N0)? mem[1021] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] : 
                         (N0)? mem[1020] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] : 
                         (N0)? mem[1019] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] : 
                         (N0)? mem[1018] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] : 
                         (N0)? mem[1017] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] : 
                         (N0)? mem[1016] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] : 
                         (N0)? mem[1015] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] : 
                         (N0)? mem[1014] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] : 
                         (N0)? mem[1013] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] : 
                         (N0)? mem[1012] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] : 
                         (N0)? mem[1011] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] : 
                         (N0)? mem[1010] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] : 
                         (N0)? mem[1009] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] : 
                         (N0)? mem[1008] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] : 
                         (N0)? mem[1007] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] : 
                         (N0)? mem[1006] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] : 
                         (N0)? mem[1005] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] : 
                         (N0)? mem[1004] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] : 
                         (N0)? mem[1003] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] : 
                         (N0)? mem[1002] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] : 
                         (N0)? mem[1001] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] : 
                         (N0)? mem[1000] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] : 
                         (N0)? mem[999] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] : 
                         (N0)? mem[998] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] : 
                         (N0)? mem[997] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] : 
                         (N0)? mem[996] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] : 
                         (N0)? mem[995] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] : 
                         (N0)? mem[994] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] : 
                         (N0)? mem[993] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] : 
                         (N0)? mem[992] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] : 
                         (N0)? mem[991] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] : 
                         (N0)? mem[990] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] : 
                         (N0)? mem[989] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] : 
                         (N0)? mem[988] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] : 
                         (N0)? mem[987] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] : 
                         (N0)? mem[986] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] : 
                         (N0)? mem[985] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] : 
                         (N0)? mem[984] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] : 
                         (N0)? mem[983] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] : 
                         (N0)? mem[982] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] : 
                         (N0)? mem[981] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] : 
                         (N0)? mem[980] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] : 
                         (N0)? mem[979] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] : 
                         (N0)? mem[978] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] : 
                         (N0)? mem[977] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] : 
                         (N0)? mem[976] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] : 
                         (N0)? mem[975] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] : 
                         (N0)? mem[974] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] : 
                         (N0)? mem[973] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] : 
                         (N0)? mem[972] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] : 
                         (N0)? mem[971] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] : 
                         (N0)? mem[970] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] : 
                         (N0)? mem[969] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] : 
                         (N0)? mem[968] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] : 
                         (N0)? mem[967] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] : 
                         (N0)? mem[966] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] : 
                         (N0)? mem[965] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] : 
                         (N0)? mem[964] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] : 
                         (N0)? mem[963] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] : 
                         (N0)? mem[962] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] : 
                         (N0)? mem[961] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] : 
                         (N0)? mem[960] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] : 
                         (N0)? mem[959] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] : 
                         (N0)? mem[958] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] : 
                         (N0)? mem[957] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] : 
                         (N0)? mem[956] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] : 
                         (N0)? mem[955] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] : 
                         (N0)? mem[954] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] : 
                         (N0)? mem[953] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] : 
                         (N0)? mem[952] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] : 
                         (N0)? mem[951] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] : 
                         (N0)? mem[950] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] : 
                         (N0)? mem[949] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] : 
                         (N0)? mem[948] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] : 
                         (N0)? mem[947] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] : 
                         (N0)? mem[946] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] : 
                         (N0)? mem[945] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] : 
                         (N0)? mem[944] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] : 
                         (N0)? mem[943] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] : 
                         (N0)? mem[942] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] : 
                         (N0)? mem[941] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] : 
                         (N0)? mem[940] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] : 
                         (N0)? mem[939] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] : 
                         (N0)? mem[938] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] : 
                         (N0)? mem[937] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] : 
                         (N0)? mem[936] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] : 
                         (N0)? mem[935] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] : 
                         (N0)? mem[934] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] : 
                         (N0)? mem[933] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] : 
                         (N0)? mem[932] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] : 
                         (N0)? mem[931] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] : 
                         (N0)? mem[930] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] : 
                         (N0)? mem[929] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] : 
                         (N0)? mem[928] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] : 
                         (N0)? mem[927] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] : 
                         (N0)? mem[926] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] : 
                         (N0)? mem[925] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] : 
                         (N0)? mem[924] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] : 
                         (N0)? mem[923] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] : 
                         (N0)? mem[922] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] : 
                         (N0)? mem[921] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] : 
                         (N0)? mem[920] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] : 
                         (N0)? mem[919] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] : 
                         (N0)? mem[918] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] : 
                         (N0)? mem[917] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] : 
                         (N0)? mem[916] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] : 
                         (N0)? mem[915] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] : 
                         (N0)? mem[914] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] : 
                         (N0)? mem[913] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] : 
                         (N0)? mem[912] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] : 
                         (N0)? mem[911] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] : 
                         (N0)? mem[910] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] : 
                         (N0)? mem[909] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] : 
                         (N0)? mem[908] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] : 
                         (N0)? mem[907] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] : 
                         (N0)? mem[906] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] : 
                         (N0)? mem[905] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] : 
                         (N0)? mem[904] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] : 
                         (N0)? mem[903] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] : 
                         (N0)? mem[902] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] : 
                         (N0)? mem[901] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] : 
                         (N0)? mem[900] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] : 
                         (N0)? mem[899] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] : 
                         (N0)? mem[898] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] : 
                         (N0)? mem[897] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] : 
                         (N0)? mem[896] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] : 
                         (N0)? mem[895] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] : 
                         (N0)? mem[894] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] : 
                         (N0)? mem[893] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] : 
                         (N0)? mem[892] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] : 
                         (N0)? mem[891] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] : 
                         (N0)? mem[890] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] : 
                         (N0)? mem[889] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] : 
                         (N0)? mem[888] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] : 
                         (N0)? mem[887] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] : 
                         (N0)? mem[886] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] : 
                         (N0)? mem[885] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] : 
                         (N0)? mem[884] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] : 
                         (N0)? mem[883] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] : 
                         (N0)? mem[882] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] : 
                         (N0)? mem[881] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] : 
                         (N0)? mem[880] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] : 
                         (N0)? mem[879] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] : 
                         (N0)? mem[878] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] : 
                         (N0)? mem[877] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] : 
                         (N0)? mem[876] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] : 
                         (N0)? mem[875] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] : 
                         (N0)? mem[874] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] : 
                         (N0)? mem[873] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] : 
                         (N0)? mem[872] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] : 
                         (N0)? mem[871] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] : 
                         (N0)? mem[870] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] : 
                         (N0)? mem[869] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] : 
                         (N0)? mem[868] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] : 
                         (N0)? mem[867] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] : 
                         (N0)? mem[866] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] : 
                         (N0)? mem[865] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] : 
                         (N0)? mem[864] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] : 
                         (N0)? mem[863] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] : 
                         (N0)? mem[862] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] : 
                         (N0)? mem[861] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] : 
                         (N0)? mem[860] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] : 
                         (N0)? mem[859] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] : 
                         (N0)? mem[858] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] : 
                         (N0)? mem[857] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] : 
                         (N0)? mem[856] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] : 
                         (N0)? mem[855] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] : 
                         (N0)? mem[854] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] : 
                         (N0)? mem[853] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] : 
                         (N0)? mem[852] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] : 
                         (N0)? mem[851] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] : 
                         (N0)? mem[850] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] : 
                         (N0)? mem[849] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] : 
                         (N0)? mem[848] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] : 
                         (N0)? mem[847] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] : 
                         (N0)? mem[846] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] : 
                         (N0)? mem[845] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] : 
                         (N0)? mem[844] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] : 
                         (N0)? mem[843] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] : 
                         (N0)? mem[842] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] : 
                         (N0)? mem[841] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] : 
                         (N0)? mem[840] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] : 
                         (N0)? mem[839] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] : 
                         (N0)? mem[838] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] : 
                         (N0)? mem[837] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] : 
                         (N0)? mem[836] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] : 
                         (N0)? mem[835] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] : 
                         (N0)? mem[834] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] : 
                         (N0)? mem[833] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] : 
                         (N0)? mem[832] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] : 
                         (N0)? mem[831] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] : 
                         (N0)? mem[830] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] : 
                         (N0)? mem[829] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] : 
                         (N0)? mem[828] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] : 
                         (N0)? mem[827] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] : 
                         (N0)? mem[826] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] : 
                         (N0)? mem[825] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] : 
                         (N0)? mem[824] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] : 
                         (N0)? mem[823] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] : 
                         (N0)? mem[822] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] : 
                         (N0)? mem[821] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] : 
                         (N0)? mem[820] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] : 
                         (N0)? mem[819] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] : 
                         (N0)? mem[818] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] : 
                         (N0)? mem[817] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] : 
                         (N0)? mem[816] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] : 
                         (N0)? mem[815] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] : 
                         (N0)? mem[814] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] : 
                         (N0)? mem[813] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] : 
                         (N0)? mem[812] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] : 
                         (N0)? mem[811] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] : 
                         (N0)? mem[810] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] : 
                         (N0)? mem[809] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] : 
                         (N0)? mem[808] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] : 
                         (N0)? mem[807] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] : 
                         (N0)? mem[806] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] : 
                         (N0)? mem[805] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] : 
                         (N0)? mem[804] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] : 
                         (N0)? mem[803] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] : 
                         (N0)? mem[802] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] : 
                         (N0)? mem[801] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] : 
                         (N0)? mem[800] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] : 
                         (N0)? mem[799] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] : 
                         (N0)? mem[798] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] : 
                         (N0)? mem[797] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] : 
                         (N0)? mem[796] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] : 
                         (N0)? mem[795] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] : 
                         (N0)? mem[794] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] : 
                         (N0)? mem[793] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] : 
                         (N0)? mem[792] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] : 
                         (N0)? mem[791] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] : 
                         (N0)? mem[790] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] : 
                         (N0)? mem[789] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] : 
                         (N0)? mem[788] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] : 
                         (N0)? mem[787] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] : 
                         (N0)? mem[786] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] : 
                         (N0)? mem[785] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] : 
                         (N0)? mem[784] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] : 
                         (N0)? mem[783] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] : 
                         (N0)? mem[782] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] : 
                         (N0)? mem[781] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] : 
                         (N0)? mem[780] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] : 
                         (N0)? mem[779] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] : 
                         (N0)? mem[778] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] : 
                         (N0)? mem[777] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] : 
                         (N0)? mem[776] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] : 
                         (N0)? mem[775] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] : 
                         (N0)? mem[774] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] : 
                         (N0)? mem[773] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] : 
                         (N0)? mem[772] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] : 
                         (N0)? mem[771] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] : 
                         (N0)? mem[770] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] : 
                         (N0)? mem[769] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] : 
                         (N0)? mem[768] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] : 
                         (N0)? mem[767] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] : 
                         (N0)? mem[766] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] : 
                         (N0)? mem[765] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] : 
                         (N0)? mem[764] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] : 
                         (N0)? mem[763] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] : 
                         (N0)? mem[762] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] : 
                         (N0)? mem[761] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] : 
                         (N0)? mem[760] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] : 
                         (N0)? mem[759] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] : 
                         (N0)? mem[758] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] : 
                         (N0)? mem[757] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] : 
                         (N0)? mem[756] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] : 
                         (N0)? mem[755] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] : 
                         (N0)? mem[754] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] : 
                         (N0)? mem[753] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] : 
                         (N0)? mem[752] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] : 
                         (N0)? mem[751] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] : 
                         (N0)? mem[750] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] : 
                         (N0)? mem[749] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] : 
                         (N0)? mem[748] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] : 
                         (N0)? mem[747] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] : 
                         (N0)? mem[746] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] : 
                         (N0)? mem[745] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] : 
                         (N0)? mem[744] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] : 
                         (N0)? mem[743] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] : 
                         (N0)? mem[742] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] : 
                         (N0)? mem[741] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] : 
                         (N0)? mem[740] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] : 
                         (N0)? mem[739] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] : 
                         (N0)? mem[738] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] : 
                         (N0)? mem[737] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] : 
                         (N0)? mem[736] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] : 
                         (N0)? mem[735] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] : 
                         (N0)? mem[734] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] : 
                         (N0)? mem[733] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] : 
                         (N0)? mem[732] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] : 
                         (N0)? mem[731] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] : 
                         (N0)? mem[730] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] : 
                         (N0)? mem[729] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] : 
                         (N0)? mem[728] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] : 
                         (N0)? mem[727] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] : 
                         (N0)? mem[726] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] : 
                         (N0)? mem[725] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] : 
                         (N0)? mem[724] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] : 
                         (N0)? mem[723] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] : 
                         (N0)? mem[722] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] : 
                         (N0)? mem[721] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] : 
                         (N0)? mem[720] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] : 
                         (N0)? mem[719] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] : 
                         (N0)? mem[718] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] : 
                         (N0)? mem[717] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] : 
                         (N0)? mem[716] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] : 
                         (N0)? mem[715] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] : 
                         (N0)? mem[714] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] : 
                         (N0)? mem[713] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] : 
                         (N0)? mem[712] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] : 
                         (N0)? mem[711] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] : 
                         (N0)? mem[710] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] : 
                         (N0)? mem[709] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] : 
                         (N0)? mem[708] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] : 
                         (N0)? mem[707] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] : 
                         (N0)? mem[706] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] : 
                         (N0)? mem[705] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] : 
                         (N0)? mem[704] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] : 
                         (N0)? mem[703] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] : 
                         (N0)? mem[702] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] : 
                         (N0)? mem[701] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] : 
                         (N0)? mem[700] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] : 
                         (N0)? mem[699] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] : 
                         (N0)? mem[698] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] : 
                         (N0)? mem[697] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] : 
                         (N0)? mem[696] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] : 
                         (N0)? mem[695] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] : 
                         (N0)? mem[694] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] : 
                         (N0)? mem[693] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] : 
                         (N0)? mem[692] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] : 
                         (N0)? mem[691] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] : 
                         (N0)? mem[690] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] : 
                         (N0)? mem[689] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] : 
                         (N0)? mem[688] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] : 
                         (N0)? mem[687] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] : 
                         (N0)? mem[686] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] : 
                         (N0)? mem[685] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] : 
                         (N0)? mem[684] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] : 
                         (N0)? mem[683] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] : 
                         (N0)? mem[682] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] : 
                         (N0)? mem[681] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] : 
                         (N0)? mem[680] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] : 
                         (N0)? mem[679] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] : 
                         (N0)? mem[678] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] : 
                         (N0)? mem[677] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] : 
                         (N0)? mem[676] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] : 
                         (N0)? mem[675] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] : 
                         (N0)? mem[674] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] : 
                         (N0)? mem[673] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] : 
                         (N0)? mem[672] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] : 
                         (N0)? mem[671] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] : 
                         (N0)? mem[670] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] : 
                         (N0)? mem[669] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] : 
                         (N0)? mem[668] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] : 
                         (N0)? mem[667] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] : 
                         (N0)? mem[666] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] : 
                         (N0)? mem[665] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] : 
                         (N0)? mem[664] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] : 
                         (N0)? mem[663] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] : 
                         (N0)? mem[662] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] : 
                         (N0)? mem[661] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] : 
                         (N0)? mem[660] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] : 
                         (N0)? mem[659] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] : 
                         (N0)? mem[658] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] : 
                         (N0)? mem[657] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] : 
                         (N0)? mem[656] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] : 
                         (N0)? mem[655] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] : 
                         (N0)? mem[654] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] : 
                         (N0)? mem[653] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] : 
                         (N0)? mem[652] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] : 
                         (N0)? mem[651] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] : 
                         (N0)? mem[650] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] : 
                         (N0)? mem[649] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] : 
                         (N0)? mem[648] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] : 
                         (N0)? mem[647] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] : 
                         (N0)? mem[646] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] : 
                         (N0)? mem[645] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] : 
                         (N0)? mem[644] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] : 
                         (N0)? mem[643] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] : 
                         (N0)? mem[642] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] : 
                         (N0)? mem[641] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] : 
                         (N0)? mem[640] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] : 
                         (N0)? mem[639] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] : 
                        (N0)? mem[638] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] : 
                        (N0)? mem[637] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] : 
                        (N0)? mem[636] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] : 
                        (N0)? mem[635] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] : 
                        (N0)? mem[634] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] : 
                        (N0)? mem[633] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] : 
                        (N0)? mem[632] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] : 
                        (N0)? mem[631] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] : 
                        (N0)? mem[630] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] : 
                        (N0)? mem[629] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] : 
                        (N0)? mem[628] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] : 
                        (N0)? mem[627] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] : 
                        (N0)? mem[626] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] : 
                        (N0)? mem[625] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] : 
                        (N0)? mem[624] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] : 
                        (N0)? mem[623] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] : 
                        (N0)? mem[622] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] : 
                        (N0)? mem[621] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] : 
                        (N0)? mem[620] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] : 
                        (N0)? mem[619] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] : 
                        (N0)? mem[618] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] : 
                        (N0)? mem[617] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] : 
                        (N0)? mem[616] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] : 
                        (N0)? mem[615] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] : 
                        (N0)? mem[614] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] : 
                        (N0)? mem[613] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] : 
                        (N0)? mem[612] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] : 
                        (N0)? mem[611] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] : 
                        (N0)? mem[610] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] : 
                        (N0)? mem[609] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] : 
                        (N0)? mem[608] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] : 
                        (N0)? mem[607] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] : 
                        (N0)? mem[606] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] : 
                        (N0)? mem[605] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] : 
                        (N0)? mem[604] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] : 
                        (N0)? mem[603] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[602] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[601] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[600] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[599] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[598] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[597] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[596] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[595] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[594] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[593] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[592] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[591] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[590] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[589] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[588] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[587] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[586] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[585] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[584] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[583] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[582] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[581] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[580] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[579] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[578] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[577] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[576] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[575] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[574] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[573] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[572] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[571] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[570] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[569] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[568] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[567] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[566] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[565] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[564] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[563] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[562] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[561] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[560] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[559] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[558] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[557] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[556] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[555] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[554] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[553] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[552] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[551] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[550] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[549] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[548] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[547] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[546] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[545] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[544] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[543] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[542] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[541] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[540] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[539] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } : 
                                                                       (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N13) begin
      { mem[1077:979], mem[539:539] } <= { w_data_i[538:440], w_data_i[0:0] };
    end 
    if(N14) begin
      { mem[978:880], mem[540:540] } <= { w_data_i[439:341], w_data_i[1:1] };
    end 
    if(N15) begin
      { mem[879:781], mem[541:541] } <= { w_data_i[340:242], w_data_i[2:2] };
    end 
    if(N16) begin
      { mem[780:682], mem[542:542] } <= { w_data_i[241:143], w_data_i[3:3] };
    end 
    if(N17) begin
      { mem[681:583], mem[543:543] } <= { w_data_i[142:44], w_data_i[4:4] };
    end 
    if(N18) begin
      { mem[582:544] } <= { w_data_i[43:5] };
    end 
    if(N7) begin
      { mem[538:440], mem[0:0] } <= { w_data_i[538:440], w_data_i[0:0] };
    end 
    if(N8) begin
      { mem[439:341], mem[1:1] } <= { w_data_i[439:341], w_data_i[1:1] };
    end 
    if(N9) begin
      { mem[340:242], mem[2:2] } <= { w_data_i[340:242], w_data_i[2:2] };
    end 
    if(N10) begin
      { mem[241:143], mem[3:3] } <= { w_data_i[241:143], w_data_i[3:3] };
    end 
    if(N11) begin
      { mem[142:44], mem[4:4] } <= { w_data_i[142:44], w_data_i[4:4] };
    end 
    if(N12) begin
      { mem[43:5] } <= { w_data_i[43:5] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p539_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [538:0] w_data_i;
  input [0:0] r_addr_i;
  output [538:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [538:0] r_data_o;

  bsg_mem_1r1w_synth_width_p539_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p539
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [538:0] data_i;
  output [538:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [538:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p539_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bp_be_dcache_lce_tr_num_lce_p2_num_cce_p1_data_width_p64_paddr_width_p22_lce_data_width_p512_ways_p8_sets_p64
(
  tr_received_o,
  lce_tr_resp_i,
  lce_tr_resp_v_i,
  lce_tr_resp_yumi_o,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_pkt_yumi_i
);

  input [538:0] lce_tr_resp_i;
  output [521:0] data_mem_pkt_o;
  input lce_tr_resp_v_i;
  input data_mem_pkt_yumi_i;
  output tr_received_o;
  output lce_tr_resp_yumi_o;
  output data_mem_pkt_v_o;
  wire [521:0] data_mem_pkt_o;
  wire tr_received_o,lce_tr_resp_yumi_o,data_mem_pkt_v_o,data_mem_pkt_yumi_i,
  lce_tr_resp_v_i;
  assign data_mem_pkt_o[0] = 1'b1;
  assign tr_received_o = data_mem_pkt_yumi_i;
  assign lce_tr_resp_yumi_o = data_mem_pkt_yumi_i;
  assign data_mem_pkt_v_o = lce_tr_resp_v_i;
  assign data_mem_pkt_o[521] = lce_tr_resp_i[523];
  assign data_mem_pkt_o[520] = lce_tr_resp_i[522];
  assign data_mem_pkt_o[519] = lce_tr_resp_i[521];
  assign data_mem_pkt_o[518] = lce_tr_resp_i[520];
  assign data_mem_pkt_o[517] = lce_tr_resp_i[519];
  assign data_mem_pkt_o[516] = lce_tr_resp_i[518];
  assign data_mem_pkt_o[515] = lce_tr_resp_i[536];
  assign data_mem_pkt_o[514] = lce_tr_resp_i[535];
  assign data_mem_pkt_o[513] = lce_tr_resp_i[534];
  assign data_mem_pkt_o[512] = lce_tr_resp_i[511];
  assign data_mem_pkt_o[511] = lce_tr_resp_i[510];
  assign data_mem_pkt_o[510] = lce_tr_resp_i[509];
  assign data_mem_pkt_o[509] = lce_tr_resp_i[508];
  assign data_mem_pkt_o[508] = lce_tr_resp_i[507];
  assign data_mem_pkt_o[507] = lce_tr_resp_i[506];
  assign data_mem_pkt_o[506] = lce_tr_resp_i[505];
  assign data_mem_pkt_o[505] = lce_tr_resp_i[504];
  assign data_mem_pkt_o[504] = lce_tr_resp_i[503];
  assign data_mem_pkt_o[503] = lce_tr_resp_i[502];
  assign data_mem_pkt_o[502] = lce_tr_resp_i[501];
  assign data_mem_pkt_o[501] = lce_tr_resp_i[500];
  assign data_mem_pkt_o[500] = lce_tr_resp_i[499];
  assign data_mem_pkt_o[499] = lce_tr_resp_i[498];
  assign data_mem_pkt_o[498] = lce_tr_resp_i[497];
  assign data_mem_pkt_o[497] = lce_tr_resp_i[496];
  assign data_mem_pkt_o[496] = lce_tr_resp_i[495];
  assign data_mem_pkt_o[495] = lce_tr_resp_i[494];
  assign data_mem_pkt_o[494] = lce_tr_resp_i[493];
  assign data_mem_pkt_o[493] = lce_tr_resp_i[492];
  assign data_mem_pkt_o[492] = lce_tr_resp_i[491];
  assign data_mem_pkt_o[491] = lce_tr_resp_i[490];
  assign data_mem_pkt_o[490] = lce_tr_resp_i[489];
  assign data_mem_pkt_o[489] = lce_tr_resp_i[488];
  assign data_mem_pkt_o[488] = lce_tr_resp_i[487];
  assign data_mem_pkt_o[487] = lce_tr_resp_i[486];
  assign data_mem_pkt_o[486] = lce_tr_resp_i[485];
  assign data_mem_pkt_o[485] = lce_tr_resp_i[484];
  assign data_mem_pkt_o[484] = lce_tr_resp_i[483];
  assign data_mem_pkt_o[483] = lce_tr_resp_i[482];
  assign data_mem_pkt_o[482] = lce_tr_resp_i[481];
  assign data_mem_pkt_o[481] = lce_tr_resp_i[480];
  assign data_mem_pkt_o[480] = lce_tr_resp_i[479];
  assign data_mem_pkt_o[479] = lce_tr_resp_i[478];
  assign data_mem_pkt_o[478] = lce_tr_resp_i[477];
  assign data_mem_pkt_o[477] = lce_tr_resp_i[476];
  assign data_mem_pkt_o[476] = lce_tr_resp_i[475];
  assign data_mem_pkt_o[475] = lce_tr_resp_i[474];
  assign data_mem_pkt_o[474] = lce_tr_resp_i[473];
  assign data_mem_pkt_o[473] = lce_tr_resp_i[472];
  assign data_mem_pkt_o[472] = lce_tr_resp_i[471];
  assign data_mem_pkt_o[471] = lce_tr_resp_i[470];
  assign data_mem_pkt_o[470] = lce_tr_resp_i[469];
  assign data_mem_pkt_o[469] = lce_tr_resp_i[468];
  assign data_mem_pkt_o[468] = lce_tr_resp_i[467];
  assign data_mem_pkt_o[467] = lce_tr_resp_i[466];
  assign data_mem_pkt_o[466] = lce_tr_resp_i[465];
  assign data_mem_pkt_o[465] = lce_tr_resp_i[464];
  assign data_mem_pkt_o[464] = lce_tr_resp_i[463];
  assign data_mem_pkt_o[463] = lce_tr_resp_i[462];
  assign data_mem_pkt_o[462] = lce_tr_resp_i[461];
  assign data_mem_pkt_o[461] = lce_tr_resp_i[460];
  assign data_mem_pkt_o[460] = lce_tr_resp_i[459];
  assign data_mem_pkt_o[459] = lce_tr_resp_i[458];
  assign data_mem_pkt_o[458] = lce_tr_resp_i[457];
  assign data_mem_pkt_o[457] = lce_tr_resp_i[456];
  assign data_mem_pkt_o[456] = lce_tr_resp_i[455];
  assign data_mem_pkt_o[455] = lce_tr_resp_i[454];
  assign data_mem_pkt_o[454] = lce_tr_resp_i[453];
  assign data_mem_pkt_o[453] = lce_tr_resp_i[452];
  assign data_mem_pkt_o[452] = lce_tr_resp_i[451];
  assign data_mem_pkt_o[451] = lce_tr_resp_i[450];
  assign data_mem_pkt_o[450] = lce_tr_resp_i[449];
  assign data_mem_pkt_o[449] = lce_tr_resp_i[448];
  assign data_mem_pkt_o[448] = lce_tr_resp_i[447];
  assign data_mem_pkt_o[447] = lce_tr_resp_i[446];
  assign data_mem_pkt_o[446] = lce_tr_resp_i[445];
  assign data_mem_pkt_o[445] = lce_tr_resp_i[444];
  assign data_mem_pkt_o[444] = lce_tr_resp_i[443];
  assign data_mem_pkt_o[443] = lce_tr_resp_i[442];
  assign data_mem_pkt_o[442] = lce_tr_resp_i[441];
  assign data_mem_pkt_o[441] = lce_tr_resp_i[440];
  assign data_mem_pkt_o[440] = lce_tr_resp_i[439];
  assign data_mem_pkt_o[439] = lce_tr_resp_i[438];
  assign data_mem_pkt_o[438] = lce_tr_resp_i[437];
  assign data_mem_pkt_o[437] = lce_tr_resp_i[436];
  assign data_mem_pkt_o[436] = lce_tr_resp_i[435];
  assign data_mem_pkt_o[435] = lce_tr_resp_i[434];
  assign data_mem_pkt_o[434] = lce_tr_resp_i[433];
  assign data_mem_pkt_o[433] = lce_tr_resp_i[432];
  assign data_mem_pkt_o[432] = lce_tr_resp_i[431];
  assign data_mem_pkt_o[431] = lce_tr_resp_i[430];
  assign data_mem_pkt_o[430] = lce_tr_resp_i[429];
  assign data_mem_pkt_o[429] = lce_tr_resp_i[428];
  assign data_mem_pkt_o[428] = lce_tr_resp_i[427];
  assign data_mem_pkt_o[427] = lce_tr_resp_i[426];
  assign data_mem_pkt_o[426] = lce_tr_resp_i[425];
  assign data_mem_pkt_o[425] = lce_tr_resp_i[424];
  assign data_mem_pkt_o[424] = lce_tr_resp_i[423];
  assign data_mem_pkt_o[423] = lce_tr_resp_i[422];
  assign data_mem_pkt_o[422] = lce_tr_resp_i[421];
  assign data_mem_pkt_o[421] = lce_tr_resp_i[420];
  assign data_mem_pkt_o[420] = lce_tr_resp_i[419];
  assign data_mem_pkt_o[419] = lce_tr_resp_i[418];
  assign data_mem_pkt_o[418] = lce_tr_resp_i[417];
  assign data_mem_pkt_o[417] = lce_tr_resp_i[416];
  assign data_mem_pkt_o[416] = lce_tr_resp_i[415];
  assign data_mem_pkt_o[415] = lce_tr_resp_i[414];
  assign data_mem_pkt_o[414] = lce_tr_resp_i[413];
  assign data_mem_pkt_o[413] = lce_tr_resp_i[412];
  assign data_mem_pkt_o[412] = lce_tr_resp_i[411];
  assign data_mem_pkt_o[411] = lce_tr_resp_i[410];
  assign data_mem_pkt_o[410] = lce_tr_resp_i[409];
  assign data_mem_pkt_o[409] = lce_tr_resp_i[408];
  assign data_mem_pkt_o[408] = lce_tr_resp_i[407];
  assign data_mem_pkt_o[407] = lce_tr_resp_i[406];
  assign data_mem_pkt_o[406] = lce_tr_resp_i[405];
  assign data_mem_pkt_o[405] = lce_tr_resp_i[404];
  assign data_mem_pkt_o[404] = lce_tr_resp_i[403];
  assign data_mem_pkt_o[403] = lce_tr_resp_i[402];
  assign data_mem_pkt_o[402] = lce_tr_resp_i[401];
  assign data_mem_pkt_o[401] = lce_tr_resp_i[400];
  assign data_mem_pkt_o[400] = lce_tr_resp_i[399];
  assign data_mem_pkt_o[399] = lce_tr_resp_i[398];
  assign data_mem_pkt_o[398] = lce_tr_resp_i[397];
  assign data_mem_pkt_o[397] = lce_tr_resp_i[396];
  assign data_mem_pkt_o[396] = lce_tr_resp_i[395];
  assign data_mem_pkt_o[395] = lce_tr_resp_i[394];
  assign data_mem_pkt_o[394] = lce_tr_resp_i[393];
  assign data_mem_pkt_o[393] = lce_tr_resp_i[392];
  assign data_mem_pkt_o[392] = lce_tr_resp_i[391];
  assign data_mem_pkt_o[391] = lce_tr_resp_i[390];
  assign data_mem_pkt_o[390] = lce_tr_resp_i[389];
  assign data_mem_pkt_o[389] = lce_tr_resp_i[388];
  assign data_mem_pkt_o[388] = lce_tr_resp_i[387];
  assign data_mem_pkt_o[387] = lce_tr_resp_i[386];
  assign data_mem_pkt_o[386] = lce_tr_resp_i[385];
  assign data_mem_pkt_o[385] = lce_tr_resp_i[384];
  assign data_mem_pkt_o[384] = lce_tr_resp_i[383];
  assign data_mem_pkt_o[383] = lce_tr_resp_i[382];
  assign data_mem_pkt_o[382] = lce_tr_resp_i[381];
  assign data_mem_pkt_o[381] = lce_tr_resp_i[380];
  assign data_mem_pkt_o[380] = lce_tr_resp_i[379];
  assign data_mem_pkt_o[379] = lce_tr_resp_i[378];
  assign data_mem_pkt_o[378] = lce_tr_resp_i[377];
  assign data_mem_pkt_o[377] = lce_tr_resp_i[376];
  assign data_mem_pkt_o[376] = lce_tr_resp_i[375];
  assign data_mem_pkt_o[375] = lce_tr_resp_i[374];
  assign data_mem_pkt_o[374] = lce_tr_resp_i[373];
  assign data_mem_pkt_o[373] = lce_tr_resp_i[372];
  assign data_mem_pkt_o[372] = lce_tr_resp_i[371];
  assign data_mem_pkt_o[371] = lce_tr_resp_i[370];
  assign data_mem_pkt_o[370] = lce_tr_resp_i[369];
  assign data_mem_pkt_o[369] = lce_tr_resp_i[368];
  assign data_mem_pkt_o[368] = lce_tr_resp_i[367];
  assign data_mem_pkt_o[367] = lce_tr_resp_i[366];
  assign data_mem_pkt_o[366] = lce_tr_resp_i[365];
  assign data_mem_pkt_o[365] = lce_tr_resp_i[364];
  assign data_mem_pkt_o[364] = lce_tr_resp_i[363];
  assign data_mem_pkt_o[363] = lce_tr_resp_i[362];
  assign data_mem_pkt_o[362] = lce_tr_resp_i[361];
  assign data_mem_pkt_o[361] = lce_tr_resp_i[360];
  assign data_mem_pkt_o[360] = lce_tr_resp_i[359];
  assign data_mem_pkt_o[359] = lce_tr_resp_i[358];
  assign data_mem_pkt_o[358] = lce_tr_resp_i[357];
  assign data_mem_pkt_o[357] = lce_tr_resp_i[356];
  assign data_mem_pkt_o[356] = lce_tr_resp_i[355];
  assign data_mem_pkt_o[355] = lce_tr_resp_i[354];
  assign data_mem_pkt_o[354] = lce_tr_resp_i[353];
  assign data_mem_pkt_o[353] = lce_tr_resp_i[352];
  assign data_mem_pkt_o[352] = lce_tr_resp_i[351];
  assign data_mem_pkt_o[351] = lce_tr_resp_i[350];
  assign data_mem_pkt_o[350] = lce_tr_resp_i[349];
  assign data_mem_pkt_o[349] = lce_tr_resp_i[348];
  assign data_mem_pkt_o[348] = lce_tr_resp_i[347];
  assign data_mem_pkt_o[347] = lce_tr_resp_i[346];
  assign data_mem_pkt_o[346] = lce_tr_resp_i[345];
  assign data_mem_pkt_o[345] = lce_tr_resp_i[344];
  assign data_mem_pkt_o[344] = lce_tr_resp_i[343];
  assign data_mem_pkt_o[343] = lce_tr_resp_i[342];
  assign data_mem_pkt_o[342] = lce_tr_resp_i[341];
  assign data_mem_pkt_o[341] = lce_tr_resp_i[340];
  assign data_mem_pkt_o[340] = lce_tr_resp_i[339];
  assign data_mem_pkt_o[339] = lce_tr_resp_i[338];
  assign data_mem_pkt_o[338] = lce_tr_resp_i[337];
  assign data_mem_pkt_o[337] = lce_tr_resp_i[336];
  assign data_mem_pkt_o[336] = lce_tr_resp_i[335];
  assign data_mem_pkt_o[335] = lce_tr_resp_i[334];
  assign data_mem_pkt_o[334] = lce_tr_resp_i[333];
  assign data_mem_pkt_o[333] = lce_tr_resp_i[332];
  assign data_mem_pkt_o[332] = lce_tr_resp_i[331];
  assign data_mem_pkt_o[331] = lce_tr_resp_i[330];
  assign data_mem_pkt_o[330] = lce_tr_resp_i[329];
  assign data_mem_pkt_o[329] = lce_tr_resp_i[328];
  assign data_mem_pkt_o[328] = lce_tr_resp_i[327];
  assign data_mem_pkt_o[327] = lce_tr_resp_i[326];
  assign data_mem_pkt_o[326] = lce_tr_resp_i[325];
  assign data_mem_pkt_o[325] = lce_tr_resp_i[324];
  assign data_mem_pkt_o[324] = lce_tr_resp_i[323];
  assign data_mem_pkt_o[323] = lce_tr_resp_i[322];
  assign data_mem_pkt_o[322] = lce_tr_resp_i[321];
  assign data_mem_pkt_o[321] = lce_tr_resp_i[320];
  assign data_mem_pkt_o[320] = lce_tr_resp_i[319];
  assign data_mem_pkt_o[319] = lce_tr_resp_i[318];
  assign data_mem_pkt_o[318] = lce_tr_resp_i[317];
  assign data_mem_pkt_o[317] = lce_tr_resp_i[316];
  assign data_mem_pkt_o[316] = lce_tr_resp_i[315];
  assign data_mem_pkt_o[315] = lce_tr_resp_i[314];
  assign data_mem_pkt_o[314] = lce_tr_resp_i[313];
  assign data_mem_pkt_o[313] = lce_tr_resp_i[312];
  assign data_mem_pkt_o[312] = lce_tr_resp_i[311];
  assign data_mem_pkt_o[311] = lce_tr_resp_i[310];
  assign data_mem_pkt_o[310] = lce_tr_resp_i[309];
  assign data_mem_pkt_o[309] = lce_tr_resp_i[308];
  assign data_mem_pkt_o[308] = lce_tr_resp_i[307];
  assign data_mem_pkt_o[307] = lce_tr_resp_i[306];
  assign data_mem_pkt_o[306] = lce_tr_resp_i[305];
  assign data_mem_pkt_o[305] = lce_tr_resp_i[304];
  assign data_mem_pkt_o[304] = lce_tr_resp_i[303];
  assign data_mem_pkt_o[303] = lce_tr_resp_i[302];
  assign data_mem_pkt_o[302] = lce_tr_resp_i[301];
  assign data_mem_pkt_o[301] = lce_tr_resp_i[300];
  assign data_mem_pkt_o[300] = lce_tr_resp_i[299];
  assign data_mem_pkt_o[299] = lce_tr_resp_i[298];
  assign data_mem_pkt_o[298] = lce_tr_resp_i[297];
  assign data_mem_pkt_o[297] = lce_tr_resp_i[296];
  assign data_mem_pkt_o[296] = lce_tr_resp_i[295];
  assign data_mem_pkt_o[295] = lce_tr_resp_i[294];
  assign data_mem_pkt_o[294] = lce_tr_resp_i[293];
  assign data_mem_pkt_o[293] = lce_tr_resp_i[292];
  assign data_mem_pkt_o[292] = lce_tr_resp_i[291];
  assign data_mem_pkt_o[291] = lce_tr_resp_i[290];
  assign data_mem_pkt_o[290] = lce_tr_resp_i[289];
  assign data_mem_pkt_o[289] = lce_tr_resp_i[288];
  assign data_mem_pkt_o[288] = lce_tr_resp_i[287];
  assign data_mem_pkt_o[287] = lce_tr_resp_i[286];
  assign data_mem_pkt_o[286] = lce_tr_resp_i[285];
  assign data_mem_pkt_o[285] = lce_tr_resp_i[284];
  assign data_mem_pkt_o[284] = lce_tr_resp_i[283];
  assign data_mem_pkt_o[283] = lce_tr_resp_i[282];
  assign data_mem_pkt_o[282] = lce_tr_resp_i[281];
  assign data_mem_pkt_o[281] = lce_tr_resp_i[280];
  assign data_mem_pkt_o[280] = lce_tr_resp_i[279];
  assign data_mem_pkt_o[279] = lce_tr_resp_i[278];
  assign data_mem_pkt_o[278] = lce_tr_resp_i[277];
  assign data_mem_pkt_o[277] = lce_tr_resp_i[276];
  assign data_mem_pkt_o[276] = lce_tr_resp_i[275];
  assign data_mem_pkt_o[275] = lce_tr_resp_i[274];
  assign data_mem_pkt_o[274] = lce_tr_resp_i[273];
  assign data_mem_pkt_o[273] = lce_tr_resp_i[272];
  assign data_mem_pkt_o[272] = lce_tr_resp_i[271];
  assign data_mem_pkt_o[271] = lce_tr_resp_i[270];
  assign data_mem_pkt_o[270] = lce_tr_resp_i[269];
  assign data_mem_pkt_o[269] = lce_tr_resp_i[268];
  assign data_mem_pkt_o[268] = lce_tr_resp_i[267];
  assign data_mem_pkt_o[267] = lce_tr_resp_i[266];
  assign data_mem_pkt_o[266] = lce_tr_resp_i[265];
  assign data_mem_pkt_o[265] = lce_tr_resp_i[264];
  assign data_mem_pkt_o[264] = lce_tr_resp_i[263];
  assign data_mem_pkt_o[263] = lce_tr_resp_i[262];
  assign data_mem_pkt_o[262] = lce_tr_resp_i[261];
  assign data_mem_pkt_o[261] = lce_tr_resp_i[260];
  assign data_mem_pkt_o[260] = lce_tr_resp_i[259];
  assign data_mem_pkt_o[259] = lce_tr_resp_i[258];
  assign data_mem_pkt_o[258] = lce_tr_resp_i[257];
  assign data_mem_pkt_o[257] = lce_tr_resp_i[256];
  assign data_mem_pkt_o[256] = lce_tr_resp_i[255];
  assign data_mem_pkt_o[255] = lce_tr_resp_i[254];
  assign data_mem_pkt_o[254] = lce_tr_resp_i[253];
  assign data_mem_pkt_o[253] = lce_tr_resp_i[252];
  assign data_mem_pkt_o[252] = lce_tr_resp_i[251];
  assign data_mem_pkt_o[251] = lce_tr_resp_i[250];
  assign data_mem_pkt_o[250] = lce_tr_resp_i[249];
  assign data_mem_pkt_o[249] = lce_tr_resp_i[248];
  assign data_mem_pkt_o[248] = lce_tr_resp_i[247];
  assign data_mem_pkt_o[247] = lce_tr_resp_i[246];
  assign data_mem_pkt_o[246] = lce_tr_resp_i[245];
  assign data_mem_pkt_o[245] = lce_tr_resp_i[244];
  assign data_mem_pkt_o[244] = lce_tr_resp_i[243];
  assign data_mem_pkt_o[243] = lce_tr_resp_i[242];
  assign data_mem_pkt_o[242] = lce_tr_resp_i[241];
  assign data_mem_pkt_o[241] = lce_tr_resp_i[240];
  assign data_mem_pkt_o[240] = lce_tr_resp_i[239];
  assign data_mem_pkt_o[239] = lce_tr_resp_i[238];
  assign data_mem_pkt_o[238] = lce_tr_resp_i[237];
  assign data_mem_pkt_o[237] = lce_tr_resp_i[236];
  assign data_mem_pkt_o[236] = lce_tr_resp_i[235];
  assign data_mem_pkt_o[235] = lce_tr_resp_i[234];
  assign data_mem_pkt_o[234] = lce_tr_resp_i[233];
  assign data_mem_pkt_o[233] = lce_tr_resp_i[232];
  assign data_mem_pkt_o[232] = lce_tr_resp_i[231];
  assign data_mem_pkt_o[231] = lce_tr_resp_i[230];
  assign data_mem_pkt_o[230] = lce_tr_resp_i[229];
  assign data_mem_pkt_o[229] = lce_tr_resp_i[228];
  assign data_mem_pkt_o[228] = lce_tr_resp_i[227];
  assign data_mem_pkt_o[227] = lce_tr_resp_i[226];
  assign data_mem_pkt_o[226] = lce_tr_resp_i[225];
  assign data_mem_pkt_o[225] = lce_tr_resp_i[224];
  assign data_mem_pkt_o[224] = lce_tr_resp_i[223];
  assign data_mem_pkt_o[223] = lce_tr_resp_i[222];
  assign data_mem_pkt_o[222] = lce_tr_resp_i[221];
  assign data_mem_pkt_o[221] = lce_tr_resp_i[220];
  assign data_mem_pkt_o[220] = lce_tr_resp_i[219];
  assign data_mem_pkt_o[219] = lce_tr_resp_i[218];
  assign data_mem_pkt_o[218] = lce_tr_resp_i[217];
  assign data_mem_pkt_o[217] = lce_tr_resp_i[216];
  assign data_mem_pkt_o[216] = lce_tr_resp_i[215];
  assign data_mem_pkt_o[215] = lce_tr_resp_i[214];
  assign data_mem_pkt_o[214] = lce_tr_resp_i[213];
  assign data_mem_pkt_o[213] = lce_tr_resp_i[212];
  assign data_mem_pkt_o[212] = lce_tr_resp_i[211];
  assign data_mem_pkt_o[211] = lce_tr_resp_i[210];
  assign data_mem_pkt_o[210] = lce_tr_resp_i[209];
  assign data_mem_pkt_o[209] = lce_tr_resp_i[208];
  assign data_mem_pkt_o[208] = lce_tr_resp_i[207];
  assign data_mem_pkt_o[207] = lce_tr_resp_i[206];
  assign data_mem_pkt_o[206] = lce_tr_resp_i[205];
  assign data_mem_pkt_o[205] = lce_tr_resp_i[204];
  assign data_mem_pkt_o[204] = lce_tr_resp_i[203];
  assign data_mem_pkt_o[203] = lce_tr_resp_i[202];
  assign data_mem_pkt_o[202] = lce_tr_resp_i[201];
  assign data_mem_pkt_o[201] = lce_tr_resp_i[200];
  assign data_mem_pkt_o[200] = lce_tr_resp_i[199];
  assign data_mem_pkt_o[199] = lce_tr_resp_i[198];
  assign data_mem_pkt_o[198] = lce_tr_resp_i[197];
  assign data_mem_pkt_o[197] = lce_tr_resp_i[196];
  assign data_mem_pkt_o[196] = lce_tr_resp_i[195];
  assign data_mem_pkt_o[195] = lce_tr_resp_i[194];
  assign data_mem_pkt_o[194] = lce_tr_resp_i[193];
  assign data_mem_pkt_o[193] = lce_tr_resp_i[192];
  assign data_mem_pkt_o[192] = lce_tr_resp_i[191];
  assign data_mem_pkt_o[191] = lce_tr_resp_i[190];
  assign data_mem_pkt_o[190] = lce_tr_resp_i[189];
  assign data_mem_pkt_o[189] = lce_tr_resp_i[188];
  assign data_mem_pkt_o[188] = lce_tr_resp_i[187];
  assign data_mem_pkt_o[187] = lce_tr_resp_i[186];
  assign data_mem_pkt_o[186] = lce_tr_resp_i[185];
  assign data_mem_pkt_o[185] = lce_tr_resp_i[184];
  assign data_mem_pkt_o[184] = lce_tr_resp_i[183];
  assign data_mem_pkt_o[183] = lce_tr_resp_i[182];
  assign data_mem_pkt_o[182] = lce_tr_resp_i[181];
  assign data_mem_pkt_o[181] = lce_tr_resp_i[180];
  assign data_mem_pkt_o[180] = lce_tr_resp_i[179];
  assign data_mem_pkt_o[179] = lce_tr_resp_i[178];
  assign data_mem_pkt_o[178] = lce_tr_resp_i[177];
  assign data_mem_pkt_o[177] = lce_tr_resp_i[176];
  assign data_mem_pkt_o[176] = lce_tr_resp_i[175];
  assign data_mem_pkt_o[175] = lce_tr_resp_i[174];
  assign data_mem_pkt_o[174] = lce_tr_resp_i[173];
  assign data_mem_pkt_o[173] = lce_tr_resp_i[172];
  assign data_mem_pkt_o[172] = lce_tr_resp_i[171];
  assign data_mem_pkt_o[171] = lce_tr_resp_i[170];
  assign data_mem_pkt_o[170] = lce_tr_resp_i[169];
  assign data_mem_pkt_o[169] = lce_tr_resp_i[168];
  assign data_mem_pkt_o[168] = lce_tr_resp_i[167];
  assign data_mem_pkt_o[167] = lce_tr_resp_i[166];
  assign data_mem_pkt_o[166] = lce_tr_resp_i[165];
  assign data_mem_pkt_o[165] = lce_tr_resp_i[164];
  assign data_mem_pkt_o[164] = lce_tr_resp_i[163];
  assign data_mem_pkt_o[163] = lce_tr_resp_i[162];
  assign data_mem_pkt_o[162] = lce_tr_resp_i[161];
  assign data_mem_pkt_o[161] = lce_tr_resp_i[160];
  assign data_mem_pkt_o[160] = lce_tr_resp_i[159];
  assign data_mem_pkt_o[159] = lce_tr_resp_i[158];
  assign data_mem_pkt_o[158] = lce_tr_resp_i[157];
  assign data_mem_pkt_o[157] = lce_tr_resp_i[156];
  assign data_mem_pkt_o[156] = lce_tr_resp_i[155];
  assign data_mem_pkt_o[155] = lce_tr_resp_i[154];
  assign data_mem_pkt_o[154] = lce_tr_resp_i[153];
  assign data_mem_pkt_o[153] = lce_tr_resp_i[152];
  assign data_mem_pkt_o[152] = lce_tr_resp_i[151];
  assign data_mem_pkt_o[151] = lce_tr_resp_i[150];
  assign data_mem_pkt_o[150] = lce_tr_resp_i[149];
  assign data_mem_pkt_o[149] = lce_tr_resp_i[148];
  assign data_mem_pkt_o[148] = lce_tr_resp_i[147];
  assign data_mem_pkt_o[147] = lce_tr_resp_i[146];
  assign data_mem_pkt_o[146] = lce_tr_resp_i[145];
  assign data_mem_pkt_o[145] = lce_tr_resp_i[144];
  assign data_mem_pkt_o[144] = lce_tr_resp_i[143];
  assign data_mem_pkt_o[143] = lce_tr_resp_i[142];
  assign data_mem_pkt_o[142] = lce_tr_resp_i[141];
  assign data_mem_pkt_o[141] = lce_tr_resp_i[140];
  assign data_mem_pkt_o[140] = lce_tr_resp_i[139];
  assign data_mem_pkt_o[139] = lce_tr_resp_i[138];
  assign data_mem_pkt_o[138] = lce_tr_resp_i[137];
  assign data_mem_pkt_o[137] = lce_tr_resp_i[136];
  assign data_mem_pkt_o[136] = lce_tr_resp_i[135];
  assign data_mem_pkt_o[135] = lce_tr_resp_i[134];
  assign data_mem_pkt_o[134] = lce_tr_resp_i[133];
  assign data_mem_pkt_o[133] = lce_tr_resp_i[132];
  assign data_mem_pkt_o[132] = lce_tr_resp_i[131];
  assign data_mem_pkt_o[131] = lce_tr_resp_i[130];
  assign data_mem_pkt_o[130] = lce_tr_resp_i[129];
  assign data_mem_pkt_o[129] = lce_tr_resp_i[128];
  assign data_mem_pkt_o[128] = lce_tr_resp_i[127];
  assign data_mem_pkt_o[127] = lce_tr_resp_i[126];
  assign data_mem_pkt_o[126] = lce_tr_resp_i[125];
  assign data_mem_pkt_o[125] = lce_tr_resp_i[124];
  assign data_mem_pkt_o[124] = lce_tr_resp_i[123];
  assign data_mem_pkt_o[123] = lce_tr_resp_i[122];
  assign data_mem_pkt_o[122] = lce_tr_resp_i[121];
  assign data_mem_pkt_o[121] = lce_tr_resp_i[120];
  assign data_mem_pkt_o[120] = lce_tr_resp_i[119];
  assign data_mem_pkt_o[119] = lce_tr_resp_i[118];
  assign data_mem_pkt_o[118] = lce_tr_resp_i[117];
  assign data_mem_pkt_o[117] = lce_tr_resp_i[116];
  assign data_mem_pkt_o[116] = lce_tr_resp_i[115];
  assign data_mem_pkt_o[115] = lce_tr_resp_i[114];
  assign data_mem_pkt_o[114] = lce_tr_resp_i[113];
  assign data_mem_pkt_o[113] = lce_tr_resp_i[112];
  assign data_mem_pkt_o[112] = lce_tr_resp_i[111];
  assign data_mem_pkt_o[111] = lce_tr_resp_i[110];
  assign data_mem_pkt_o[110] = lce_tr_resp_i[109];
  assign data_mem_pkt_o[109] = lce_tr_resp_i[108];
  assign data_mem_pkt_o[108] = lce_tr_resp_i[107];
  assign data_mem_pkt_o[107] = lce_tr_resp_i[106];
  assign data_mem_pkt_o[106] = lce_tr_resp_i[105];
  assign data_mem_pkt_o[105] = lce_tr_resp_i[104];
  assign data_mem_pkt_o[104] = lce_tr_resp_i[103];
  assign data_mem_pkt_o[103] = lce_tr_resp_i[102];
  assign data_mem_pkt_o[102] = lce_tr_resp_i[101];
  assign data_mem_pkt_o[101] = lce_tr_resp_i[100];
  assign data_mem_pkt_o[100] = lce_tr_resp_i[99];
  assign data_mem_pkt_o[99] = lce_tr_resp_i[98];
  assign data_mem_pkt_o[98] = lce_tr_resp_i[97];
  assign data_mem_pkt_o[97] = lce_tr_resp_i[96];
  assign data_mem_pkt_o[96] = lce_tr_resp_i[95];
  assign data_mem_pkt_o[95] = lce_tr_resp_i[94];
  assign data_mem_pkt_o[94] = lce_tr_resp_i[93];
  assign data_mem_pkt_o[93] = lce_tr_resp_i[92];
  assign data_mem_pkt_o[92] = lce_tr_resp_i[91];
  assign data_mem_pkt_o[91] = lce_tr_resp_i[90];
  assign data_mem_pkt_o[90] = lce_tr_resp_i[89];
  assign data_mem_pkt_o[89] = lce_tr_resp_i[88];
  assign data_mem_pkt_o[88] = lce_tr_resp_i[87];
  assign data_mem_pkt_o[87] = lce_tr_resp_i[86];
  assign data_mem_pkt_o[86] = lce_tr_resp_i[85];
  assign data_mem_pkt_o[85] = lce_tr_resp_i[84];
  assign data_mem_pkt_o[84] = lce_tr_resp_i[83];
  assign data_mem_pkt_o[83] = lce_tr_resp_i[82];
  assign data_mem_pkt_o[82] = lce_tr_resp_i[81];
  assign data_mem_pkt_o[81] = lce_tr_resp_i[80];
  assign data_mem_pkt_o[80] = lce_tr_resp_i[79];
  assign data_mem_pkt_o[79] = lce_tr_resp_i[78];
  assign data_mem_pkt_o[78] = lce_tr_resp_i[77];
  assign data_mem_pkt_o[77] = lce_tr_resp_i[76];
  assign data_mem_pkt_o[76] = lce_tr_resp_i[75];
  assign data_mem_pkt_o[75] = lce_tr_resp_i[74];
  assign data_mem_pkt_o[74] = lce_tr_resp_i[73];
  assign data_mem_pkt_o[73] = lce_tr_resp_i[72];
  assign data_mem_pkt_o[72] = lce_tr_resp_i[71];
  assign data_mem_pkt_o[71] = lce_tr_resp_i[70];
  assign data_mem_pkt_o[70] = lce_tr_resp_i[69];
  assign data_mem_pkt_o[69] = lce_tr_resp_i[68];
  assign data_mem_pkt_o[68] = lce_tr_resp_i[67];
  assign data_mem_pkt_o[67] = lce_tr_resp_i[66];
  assign data_mem_pkt_o[66] = lce_tr_resp_i[65];
  assign data_mem_pkt_o[65] = lce_tr_resp_i[64];
  assign data_mem_pkt_o[64] = lce_tr_resp_i[63];
  assign data_mem_pkt_o[63] = lce_tr_resp_i[62];
  assign data_mem_pkt_o[62] = lce_tr_resp_i[61];
  assign data_mem_pkt_o[61] = lce_tr_resp_i[60];
  assign data_mem_pkt_o[60] = lce_tr_resp_i[59];
  assign data_mem_pkt_o[59] = lce_tr_resp_i[58];
  assign data_mem_pkt_o[58] = lce_tr_resp_i[57];
  assign data_mem_pkt_o[57] = lce_tr_resp_i[56];
  assign data_mem_pkt_o[56] = lce_tr_resp_i[55];
  assign data_mem_pkt_o[55] = lce_tr_resp_i[54];
  assign data_mem_pkt_o[54] = lce_tr_resp_i[53];
  assign data_mem_pkt_o[53] = lce_tr_resp_i[52];
  assign data_mem_pkt_o[52] = lce_tr_resp_i[51];
  assign data_mem_pkt_o[51] = lce_tr_resp_i[50];
  assign data_mem_pkt_o[50] = lce_tr_resp_i[49];
  assign data_mem_pkt_o[49] = lce_tr_resp_i[48];
  assign data_mem_pkt_o[48] = lce_tr_resp_i[47];
  assign data_mem_pkt_o[47] = lce_tr_resp_i[46];
  assign data_mem_pkt_o[46] = lce_tr_resp_i[45];
  assign data_mem_pkt_o[45] = lce_tr_resp_i[44];
  assign data_mem_pkt_o[44] = lce_tr_resp_i[43];
  assign data_mem_pkt_o[43] = lce_tr_resp_i[42];
  assign data_mem_pkt_o[42] = lce_tr_resp_i[41];
  assign data_mem_pkt_o[41] = lce_tr_resp_i[40];
  assign data_mem_pkt_o[40] = lce_tr_resp_i[39];
  assign data_mem_pkt_o[39] = lce_tr_resp_i[38];
  assign data_mem_pkt_o[38] = lce_tr_resp_i[37];
  assign data_mem_pkt_o[37] = lce_tr_resp_i[36];
  assign data_mem_pkt_o[36] = lce_tr_resp_i[35];
  assign data_mem_pkt_o[35] = lce_tr_resp_i[34];
  assign data_mem_pkt_o[34] = lce_tr_resp_i[33];
  assign data_mem_pkt_o[33] = lce_tr_resp_i[32];
  assign data_mem_pkt_o[32] = lce_tr_resp_i[31];
  assign data_mem_pkt_o[31] = lce_tr_resp_i[30];
  assign data_mem_pkt_o[30] = lce_tr_resp_i[29];
  assign data_mem_pkt_o[29] = lce_tr_resp_i[28];
  assign data_mem_pkt_o[28] = lce_tr_resp_i[27];
  assign data_mem_pkt_o[27] = lce_tr_resp_i[26];
  assign data_mem_pkt_o[26] = lce_tr_resp_i[25];
  assign data_mem_pkt_o[25] = lce_tr_resp_i[24];
  assign data_mem_pkt_o[24] = lce_tr_resp_i[23];
  assign data_mem_pkt_o[23] = lce_tr_resp_i[22];
  assign data_mem_pkt_o[22] = lce_tr_resp_i[21];
  assign data_mem_pkt_o[21] = lce_tr_resp_i[20];
  assign data_mem_pkt_o[20] = lce_tr_resp_i[19];
  assign data_mem_pkt_o[19] = lce_tr_resp_i[18];
  assign data_mem_pkt_o[18] = lce_tr_resp_i[17];
  assign data_mem_pkt_o[17] = lce_tr_resp_i[16];
  assign data_mem_pkt_o[16] = lce_tr_resp_i[15];
  assign data_mem_pkt_o[15] = lce_tr_resp_i[14];
  assign data_mem_pkt_o[14] = lce_tr_resp_i[13];
  assign data_mem_pkt_o[13] = lce_tr_resp_i[12];
  assign data_mem_pkt_o[12] = lce_tr_resp_i[11];
  assign data_mem_pkt_o[11] = lce_tr_resp_i[10];
  assign data_mem_pkt_o[10] = lce_tr_resp_i[9];
  assign data_mem_pkt_o[9] = lce_tr_resp_i[8];
  assign data_mem_pkt_o[8] = lce_tr_resp_i[7];
  assign data_mem_pkt_o[7] = lce_tr_resp_i[6];
  assign data_mem_pkt_o[6] = lce_tr_resp_i[5];
  assign data_mem_pkt_o[5] = lce_tr_resp_i[4];
  assign data_mem_pkt_o[4] = lce_tr_resp_i[3];
  assign data_mem_pkt_o[3] = lce_tr_resp_i[2];
  assign data_mem_pkt_o[2] = lce_tr_resp_i[1];
  assign data_mem_pkt_o[1] = lce_tr_resp_i[0];

endmodule



module bp_be_dcache_lce_data_width_p64_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_num_cce_p1_num_lce_p2
(
  clk_i,
  reset_i,
  lce_id_i,
  ready_o,
  cache_miss_o,
  load_miss_i,
  store_miss_i,
  miss_addr_i,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_data_i,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_v_o,
  tag_mem_pkt_o,
  tag_mem_pkt_yumi_i,
  stat_mem_pkt_v_o,
  stat_mem_pkt_o,
  lru_way_i,
  dirty_i,
  stat_mem_pkt_yumi_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_tr_resp_i,
  lce_tr_resp_v_i,
  lce_tr_resp_ready_o,
  lce_tr_resp_o,
  lce_tr_resp_v_o,
  lce_tr_resp_ready_i
);

  input [0:0] lce_id_i;
  input [21:0] miss_addr_i;
  output [521:0] data_mem_pkt_o;
  input [511:0] data_mem_data_i;
  output [22:0] tag_mem_pkt_o;
  output [10:0] stat_mem_pkt_o;
  input [2:0] lru_way_i;
  input [7:0] dirty_i;
  output [29:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [539:0] lce_data_cmd_i;
  input [538:0] lce_tr_resp_i;
  output [538:0] lce_tr_resp_o;
  input clk_i;
  input reset_i;
  input load_miss_i;
  input store_miss_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input stat_mem_pkt_yumi_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_tr_resp_v_i;
  input lce_tr_resp_ready_i;
  output ready_o;
  output cache_miss_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output stat_mem_pkt_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_tr_resp_ready_o;
  output lce_tr_resp_v_o;
  wire [521:0] data_mem_pkt_o,lce_cmd_data_mem_pkt_lo,lce_data_cmd_data_mem_pkt_lo,
  lce_tr_resp_in_data_mem_pkt_lo;
  wire [22:0] tag_mem_pkt_o;
  wire [10:0] stat_mem_pkt_o;
  wire [29:0] lce_req_o;
  wire [25:0] lce_resp_o,lce_req_to_lce_resp_lo,lce_cmd_to_lce_resp_lo;
  wire [536:0] lce_data_resp_o;
  wire [538:0] lce_tr_resp_o,lce_tr_resp_in_fifo_data_lo;
  wire ready_o,cache_miss_o,data_mem_pkt_v_o,tag_mem_pkt_v_o,stat_mem_pkt_v_o,
  lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,lce_data_cmd_ready_o,
  lce_tr_resp_ready_o,lce_tr_resp_v_o,N0,N1,N2,N3,N4,N5,N6,tr_received_li,
  cce_data_received_li,tag_set_li,tag_set_wakeup_li,lce_req_to_lce_resp_v_lo,
  lce_req_to_lce_resp_yumi_li,lce_cmd_fifo_v_lo,lce_cmd_fifo_yumi_li,lce_sync_done_lo,
  lce_cmd_to_lce_resp_v_lo,lce_cmd_to_lce_resp_yumi_li,lce_cmd_data_mem_pkt_v_lo,
  lce_cmd_data_mem_pkt_yumi_li,lce_data_cmd_fifo_v_lo,lce_data_cmd_fifo_yumi_li,
  lce_data_cmd_data_mem_pkt_v_lo,lce_data_cmd_data_mem_pkt_yumi_li,lce_tr_resp_in_fifo_v_lo,
  lce_tr_resp_in_fifo_yumi_li,lce_tr_resp_in_data_mem_pkt_v_lo,
  lce_tr_resp_in_data_mem_pkt_yumi_li,N7,N8,N9,N10,N11,N12,N13,timeout,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,
  N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40;
  wire [35:0] lce_cmd_fifo_data_lo;
  wire [539:0] lce_data_cmd_fifo_data_lo;
  wire [2:0] timeout_count_n;
  reg [2:0] timeout_count_r;

  bp_be_dcache_lce_req_data_width_p64_paddr_width_p22_num_cce_p1_num_lce_p2_ways_p8_sets_p64
  lce_cce_req_inst
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_id_i(lce_id_i[0]),
    .load_miss_i(load_miss_i),
    .store_miss_i(store_miss_i),
    .miss_addr_i(miss_addr_i),
    .lru_way_i(lru_way_i),
    .dirty_i(dirty_i),
    .cache_miss_o(cache_miss_o),
    .tr_received_i(tr_received_li),
    .cce_data_received_i(cce_data_received_li),
    .tag_set_i(tag_set_li),
    .tag_set_wakeup_i(tag_set_wakeup_li),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_req_to_lce_resp_lo),
    .lce_resp_v_o(lce_req_to_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_req_to_lce_resp_yumi_li)
  );


  bsg_two_fifo_width_p36
  lce_cmd_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_cmd_ready_o),
    .data_i(lce_cmd_i),
    .v_i(lce_cmd_v_i),
    .v_o(lce_cmd_fifo_v_lo),
    .data_o(lce_cmd_fifo_data_lo),
    .yumi_i(lce_cmd_fifo_yumi_li)
  );


  bp_be_dcache_lce_cmd_num_cce_p1_num_lce_p2_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_data_width_p64
  lce_cmd_inst
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_id_i(lce_id_i[0]),
    .lce_sync_done_o(lce_sync_done_lo),
    .tag_set_o(tag_set_li),
    .tag_set_wakeup_o(tag_set_wakeup_li),
    .lce_cmd_i(lce_cmd_fifo_data_lo),
    .lce_cmd_v_i(lce_cmd_fifo_v_lo),
    .lce_cmd_yumi_o(lce_cmd_fifo_yumi_li),
    .lce_resp_o(lce_cmd_to_lce_resp_lo),
    .lce_resp_v_o(lce_cmd_to_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_cmd_to_lce_resp_yumi_li),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_tr_resp_o(lce_tr_resp_o),
    .lce_tr_resp_v_o(lce_tr_resp_v_o),
    .lce_tr_resp_ready_i(lce_tr_resp_ready_i),
    .data_mem_pkt_v_o(lce_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_cmd_data_mem_pkt_lo),
    .data_mem_data_i(data_mem_data_i),
    .data_mem_pkt_yumi_i(lce_cmd_data_mem_pkt_yumi_li),
    .tag_mem_pkt_v_o(tag_mem_pkt_v_o),
    .tag_mem_pkt_o(tag_mem_pkt_o),
    .tag_mem_pkt_yumi_i(tag_mem_pkt_yumi_i),
    .stat_mem_pkt_v_o(stat_mem_pkt_v_o),
    .stat_mem_pkt_o(stat_mem_pkt_o),
    .dirty_i(dirty_i),
    .stat_mem_pkt_yumi_i(stat_mem_pkt_yumi_i)
  );


  bsg_two_fifo_width_p540
  lce_data_cmd_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_data_cmd_ready_o),
    .data_i(lce_data_cmd_i),
    .v_i(lce_data_cmd_v_i),
    .v_o(lce_data_cmd_fifo_v_lo),
    .data_o(lce_data_cmd_fifo_data_lo),
    .yumi_i(lce_data_cmd_fifo_yumi_li)
  );


  bp_be_dcache_lce_data_cmd_num_cce_p1_num_lce_p2_data_width_p64_paddr_width_p22_lce_data_width_p512_ways_p8_sets_p64
  lce_data_cmd_inst
  (
    .cce_data_received_o(cce_data_received_li),
    .lce_data_cmd_i(lce_data_cmd_fifo_data_lo),
    .lce_data_cmd_v_i(lce_data_cmd_fifo_v_lo),
    .lce_data_cmd_yumi_o(lce_data_cmd_fifo_yumi_li),
    .data_mem_pkt_v_o(lce_data_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_data_cmd_data_mem_pkt_lo),
    .data_mem_pkt_yumi_i(lce_data_cmd_data_mem_pkt_yumi_li)
  );


  bsg_two_fifo_width_p539
  lce_tr_resp_in_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_tr_resp_ready_o),
    .data_i(lce_tr_resp_i),
    .v_i(lce_tr_resp_v_i),
    .v_o(lce_tr_resp_in_fifo_v_lo),
    .data_o(lce_tr_resp_in_fifo_data_lo),
    .yumi_i(lce_tr_resp_in_fifo_yumi_li)
  );


  bp_be_dcache_lce_tr_num_lce_p2_num_cce_p1_data_width_p64_paddr_width_p22_lce_data_width_p512_ways_p8_sets_p64
  lce_tr_inst
  (
    .tr_received_o(tr_received_li),
    .lce_tr_resp_i(lce_tr_resp_in_fifo_data_lo),
    .lce_tr_resp_v_i(lce_tr_resp_in_fifo_v_lo),
    .lce_tr_resp_yumi_o(lce_tr_resp_in_fifo_yumi_li),
    .data_mem_pkt_v_o(lce_tr_resp_in_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_tr_resp_in_data_mem_pkt_lo),
    .data_mem_pkt_yumi_i(lce_tr_resp_in_data_mem_pkt_yumi_li)
  );

  assign N29 = ~timeout_count_r[2];
  assign N30 = timeout_count_r[1] | N29;
  assign N31 = timeout_count_r[0] | N30;
  assign N32 = ~N31;
  assign { N22, N21, N20 } = timeout_count_r + 1'b1;
  assign data_mem_pkt_v_o = (N0)? 1'b1 : 
                            (N10)? 1'b1 : 
                            (N8)? lce_cmd_data_mem_pkt_v_lo : 1'b0;
  assign N0 = lce_tr_resp_in_data_mem_pkt_v_lo;
  assign data_mem_pkt_o = (N0)? lce_tr_resp_in_data_mem_pkt_lo : 
                          (N10)? lce_data_cmd_data_mem_pkt_lo : 
                          (N8)? lce_cmd_data_mem_pkt_lo : 1'b0;
  assign lce_tr_resp_in_data_mem_pkt_yumi_li = (N0)? data_mem_pkt_yumi_i : 
                                               (N9)? 1'b0 : 
                                               (N1)? 1'b0 : 1'b0;
  assign N1 = 1'b0;
  assign lce_data_cmd_data_mem_pkt_yumi_li = (N0)? 1'b0 : 
                                             (N10)? data_mem_pkt_yumi_i : 
                                             (N8)? 1'b0 : 1'b0;
  assign lce_cmd_data_mem_pkt_yumi_li = (N0)? 1'b0 : 
                                        (N10)? 1'b0 : 
                                        (N8)? data_mem_pkt_yumi_i : 1'b0;
  assign lce_resp_v_o = (N2)? 1'b1 : 
                        (N3)? lce_cmd_to_lce_resp_v_lo : 1'b0;
  assign N2 = lce_req_to_lce_resp_v_lo;
  assign N3 = N11;
  assign lce_resp_o = (N2)? lce_req_to_lce_resp_lo : 
                      (N3)? lce_cmd_to_lce_resp_lo : 1'b0;
  assign lce_req_to_lce_resp_yumi_li = (N2)? lce_resp_ready_i : 
                                       (N3)? 1'b0 : 1'b0;
  assign lce_cmd_to_lce_resp_yumi_li = (N2)? 1'b0 : 
                                       (N3)? N12 : 1'b0;
  assign { N25, N24, N23 } = (N4)? { N22, N21, N20 } : 
                             (N19)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = N18;
  assign { N28, N27, N26 } = (N5)? { N25, N24, N23 } : 
                             (N16)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N15;
  assign timeout_count_n = (N6)? { 1'b0, 1'b0, 1'b0 } : 
                           (N13)? { N28, N27, N26 } : 1'b0;
  assign N6 = timeout;
  assign N7 = lce_data_cmd_data_mem_pkt_v_lo | lce_tr_resp_in_data_mem_pkt_v_lo;
  assign N8 = ~N7;
  assign N9 = ~lce_tr_resp_in_data_mem_pkt_v_lo;
  assign N10 = lce_data_cmd_data_mem_pkt_v_lo & N9;
  assign N11 = ~lce_req_to_lce_resp_v_lo;
  assign N12 = lce_cmd_to_lce_resp_v_lo & lce_resp_ready_i;
  assign timeout = N32;
  assign N13 = ~timeout;
  assign N14 = N13;
  assign N15 = N33 | stat_mem_pkt_v_o;
  assign N33 = data_mem_pkt_v_o | tag_mem_pkt_v_o;
  assign N16 = ~N15;
  assign N17 = N14 & N15;
  assign N18 = N36 & N37;
  assign N36 = N34 & N35;
  assign N34 = ~data_mem_pkt_yumi_i;
  assign N35 = ~tag_mem_pkt_yumi_i;
  assign N37 = ~stat_mem_pkt_yumi_i;
  assign N19 = ~N18;
  assign ready_o = N39 & N40;
  assign N39 = lce_sync_done_lo & N38;
  assign N38 = ~timeout;
  assign N40 = ~cache_miss_o;

  always @(posedge clk_i) begin
    if(reset_i) begin
      { timeout_count_r[2:0] } <= { 1'b0, 1'b0, 1'b0 };
    end else if(1'b1) begin
      { timeout_count_r[2:0] } <= { timeout_count_n[2:0] };
    end 
  end


endmodule



module bsg_mux_width_p64_els_p8
(
  data_i,
  sel_i,
  data_o
);

  input [511:0] data_i;
  input [2:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  assign data_o[63] = (N7)? data_i[63] : 
                      (N9)? data_i[127] : 
                      (N11)? data_i[191] : 
                      (N13)? data_i[255] : 
                      (N8)? data_i[319] : 
                      (N10)? data_i[383] : 
                      (N12)? data_i[447] : 
                      (N14)? data_i[511] : 1'b0;
  assign data_o[62] = (N7)? data_i[62] : 
                      (N9)? data_i[126] : 
                      (N11)? data_i[190] : 
                      (N13)? data_i[254] : 
                      (N8)? data_i[318] : 
                      (N10)? data_i[382] : 
                      (N12)? data_i[446] : 
                      (N14)? data_i[510] : 1'b0;
  assign data_o[61] = (N7)? data_i[61] : 
                      (N9)? data_i[125] : 
                      (N11)? data_i[189] : 
                      (N13)? data_i[253] : 
                      (N8)? data_i[317] : 
                      (N10)? data_i[381] : 
                      (N12)? data_i[445] : 
                      (N14)? data_i[509] : 1'b0;
  assign data_o[60] = (N7)? data_i[60] : 
                      (N9)? data_i[124] : 
                      (N11)? data_i[188] : 
                      (N13)? data_i[252] : 
                      (N8)? data_i[316] : 
                      (N10)? data_i[380] : 
                      (N12)? data_i[444] : 
                      (N14)? data_i[508] : 1'b0;
  assign data_o[59] = (N7)? data_i[59] : 
                      (N9)? data_i[123] : 
                      (N11)? data_i[187] : 
                      (N13)? data_i[251] : 
                      (N8)? data_i[315] : 
                      (N10)? data_i[379] : 
                      (N12)? data_i[443] : 
                      (N14)? data_i[507] : 1'b0;
  assign data_o[58] = (N7)? data_i[58] : 
                      (N9)? data_i[122] : 
                      (N11)? data_i[186] : 
                      (N13)? data_i[250] : 
                      (N8)? data_i[314] : 
                      (N10)? data_i[378] : 
                      (N12)? data_i[442] : 
                      (N14)? data_i[506] : 1'b0;
  assign data_o[57] = (N7)? data_i[57] : 
                      (N9)? data_i[121] : 
                      (N11)? data_i[185] : 
                      (N13)? data_i[249] : 
                      (N8)? data_i[313] : 
                      (N10)? data_i[377] : 
                      (N12)? data_i[441] : 
                      (N14)? data_i[505] : 1'b0;
  assign data_o[56] = (N7)? data_i[56] : 
                      (N9)? data_i[120] : 
                      (N11)? data_i[184] : 
                      (N13)? data_i[248] : 
                      (N8)? data_i[312] : 
                      (N10)? data_i[376] : 
                      (N12)? data_i[440] : 
                      (N14)? data_i[504] : 1'b0;
  assign data_o[55] = (N7)? data_i[55] : 
                      (N9)? data_i[119] : 
                      (N11)? data_i[183] : 
                      (N13)? data_i[247] : 
                      (N8)? data_i[311] : 
                      (N10)? data_i[375] : 
                      (N12)? data_i[439] : 
                      (N14)? data_i[503] : 1'b0;
  assign data_o[54] = (N7)? data_i[54] : 
                      (N9)? data_i[118] : 
                      (N11)? data_i[182] : 
                      (N13)? data_i[246] : 
                      (N8)? data_i[310] : 
                      (N10)? data_i[374] : 
                      (N12)? data_i[438] : 
                      (N14)? data_i[502] : 1'b0;
  assign data_o[53] = (N7)? data_i[53] : 
                      (N9)? data_i[117] : 
                      (N11)? data_i[181] : 
                      (N13)? data_i[245] : 
                      (N8)? data_i[309] : 
                      (N10)? data_i[373] : 
                      (N12)? data_i[437] : 
                      (N14)? data_i[501] : 1'b0;
  assign data_o[52] = (N7)? data_i[52] : 
                      (N9)? data_i[116] : 
                      (N11)? data_i[180] : 
                      (N13)? data_i[244] : 
                      (N8)? data_i[308] : 
                      (N10)? data_i[372] : 
                      (N12)? data_i[436] : 
                      (N14)? data_i[500] : 1'b0;
  assign data_o[51] = (N7)? data_i[51] : 
                      (N9)? data_i[115] : 
                      (N11)? data_i[179] : 
                      (N13)? data_i[243] : 
                      (N8)? data_i[307] : 
                      (N10)? data_i[371] : 
                      (N12)? data_i[435] : 
                      (N14)? data_i[499] : 1'b0;
  assign data_o[50] = (N7)? data_i[50] : 
                      (N9)? data_i[114] : 
                      (N11)? data_i[178] : 
                      (N13)? data_i[242] : 
                      (N8)? data_i[306] : 
                      (N10)? data_i[370] : 
                      (N12)? data_i[434] : 
                      (N14)? data_i[498] : 1'b0;
  assign data_o[49] = (N7)? data_i[49] : 
                      (N9)? data_i[113] : 
                      (N11)? data_i[177] : 
                      (N13)? data_i[241] : 
                      (N8)? data_i[305] : 
                      (N10)? data_i[369] : 
                      (N12)? data_i[433] : 
                      (N14)? data_i[497] : 1'b0;
  assign data_o[48] = (N7)? data_i[48] : 
                      (N9)? data_i[112] : 
                      (N11)? data_i[176] : 
                      (N13)? data_i[240] : 
                      (N8)? data_i[304] : 
                      (N10)? data_i[368] : 
                      (N12)? data_i[432] : 
                      (N14)? data_i[496] : 1'b0;
  assign data_o[47] = (N7)? data_i[47] : 
                      (N9)? data_i[111] : 
                      (N11)? data_i[175] : 
                      (N13)? data_i[239] : 
                      (N8)? data_i[303] : 
                      (N10)? data_i[367] : 
                      (N12)? data_i[431] : 
                      (N14)? data_i[495] : 1'b0;
  assign data_o[46] = (N7)? data_i[46] : 
                      (N9)? data_i[110] : 
                      (N11)? data_i[174] : 
                      (N13)? data_i[238] : 
                      (N8)? data_i[302] : 
                      (N10)? data_i[366] : 
                      (N12)? data_i[430] : 
                      (N14)? data_i[494] : 1'b0;
  assign data_o[45] = (N7)? data_i[45] : 
                      (N9)? data_i[109] : 
                      (N11)? data_i[173] : 
                      (N13)? data_i[237] : 
                      (N8)? data_i[301] : 
                      (N10)? data_i[365] : 
                      (N12)? data_i[429] : 
                      (N14)? data_i[493] : 1'b0;
  assign data_o[44] = (N7)? data_i[44] : 
                      (N9)? data_i[108] : 
                      (N11)? data_i[172] : 
                      (N13)? data_i[236] : 
                      (N8)? data_i[300] : 
                      (N10)? data_i[364] : 
                      (N12)? data_i[428] : 
                      (N14)? data_i[492] : 1'b0;
  assign data_o[43] = (N7)? data_i[43] : 
                      (N9)? data_i[107] : 
                      (N11)? data_i[171] : 
                      (N13)? data_i[235] : 
                      (N8)? data_i[299] : 
                      (N10)? data_i[363] : 
                      (N12)? data_i[427] : 
                      (N14)? data_i[491] : 1'b0;
  assign data_o[42] = (N7)? data_i[42] : 
                      (N9)? data_i[106] : 
                      (N11)? data_i[170] : 
                      (N13)? data_i[234] : 
                      (N8)? data_i[298] : 
                      (N10)? data_i[362] : 
                      (N12)? data_i[426] : 
                      (N14)? data_i[490] : 1'b0;
  assign data_o[41] = (N7)? data_i[41] : 
                      (N9)? data_i[105] : 
                      (N11)? data_i[169] : 
                      (N13)? data_i[233] : 
                      (N8)? data_i[297] : 
                      (N10)? data_i[361] : 
                      (N12)? data_i[425] : 
                      (N14)? data_i[489] : 1'b0;
  assign data_o[40] = (N7)? data_i[40] : 
                      (N9)? data_i[104] : 
                      (N11)? data_i[168] : 
                      (N13)? data_i[232] : 
                      (N8)? data_i[296] : 
                      (N10)? data_i[360] : 
                      (N12)? data_i[424] : 
                      (N14)? data_i[488] : 1'b0;
  assign data_o[39] = (N7)? data_i[39] : 
                      (N9)? data_i[103] : 
                      (N11)? data_i[167] : 
                      (N13)? data_i[231] : 
                      (N8)? data_i[295] : 
                      (N10)? data_i[359] : 
                      (N12)? data_i[423] : 
                      (N14)? data_i[487] : 1'b0;
  assign data_o[38] = (N7)? data_i[38] : 
                      (N9)? data_i[102] : 
                      (N11)? data_i[166] : 
                      (N13)? data_i[230] : 
                      (N8)? data_i[294] : 
                      (N10)? data_i[358] : 
                      (N12)? data_i[422] : 
                      (N14)? data_i[486] : 1'b0;
  assign data_o[37] = (N7)? data_i[37] : 
                      (N9)? data_i[101] : 
                      (N11)? data_i[165] : 
                      (N13)? data_i[229] : 
                      (N8)? data_i[293] : 
                      (N10)? data_i[357] : 
                      (N12)? data_i[421] : 
                      (N14)? data_i[485] : 1'b0;
  assign data_o[36] = (N7)? data_i[36] : 
                      (N9)? data_i[100] : 
                      (N11)? data_i[164] : 
                      (N13)? data_i[228] : 
                      (N8)? data_i[292] : 
                      (N10)? data_i[356] : 
                      (N12)? data_i[420] : 
                      (N14)? data_i[484] : 1'b0;
  assign data_o[35] = (N7)? data_i[35] : 
                      (N9)? data_i[99] : 
                      (N11)? data_i[163] : 
                      (N13)? data_i[227] : 
                      (N8)? data_i[291] : 
                      (N10)? data_i[355] : 
                      (N12)? data_i[419] : 
                      (N14)? data_i[483] : 1'b0;
  assign data_o[34] = (N7)? data_i[34] : 
                      (N9)? data_i[98] : 
                      (N11)? data_i[162] : 
                      (N13)? data_i[226] : 
                      (N8)? data_i[290] : 
                      (N10)? data_i[354] : 
                      (N12)? data_i[418] : 
                      (N14)? data_i[482] : 1'b0;
  assign data_o[33] = (N7)? data_i[33] : 
                      (N9)? data_i[97] : 
                      (N11)? data_i[161] : 
                      (N13)? data_i[225] : 
                      (N8)? data_i[289] : 
                      (N10)? data_i[353] : 
                      (N12)? data_i[417] : 
                      (N14)? data_i[481] : 1'b0;
  assign data_o[32] = (N7)? data_i[32] : 
                      (N9)? data_i[96] : 
                      (N11)? data_i[160] : 
                      (N13)? data_i[224] : 
                      (N8)? data_i[288] : 
                      (N10)? data_i[352] : 
                      (N12)? data_i[416] : 
                      (N14)? data_i[480] : 1'b0;
  assign data_o[31] = (N7)? data_i[31] : 
                      (N9)? data_i[95] : 
                      (N11)? data_i[159] : 
                      (N13)? data_i[223] : 
                      (N8)? data_i[287] : 
                      (N10)? data_i[351] : 
                      (N12)? data_i[415] : 
                      (N14)? data_i[479] : 1'b0;
  assign data_o[30] = (N7)? data_i[30] : 
                      (N9)? data_i[94] : 
                      (N11)? data_i[158] : 
                      (N13)? data_i[222] : 
                      (N8)? data_i[286] : 
                      (N10)? data_i[350] : 
                      (N12)? data_i[414] : 
                      (N14)? data_i[478] : 1'b0;
  assign data_o[29] = (N7)? data_i[29] : 
                      (N9)? data_i[93] : 
                      (N11)? data_i[157] : 
                      (N13)? data_i[221] : 
                      (N8)? data_i[285] : 
                      (N10)? data_i[349] : 
                      (N12)? data_i[413] : 
                      (N14)? data_i[477] : 1'b0;
  assign data_o[28] = (N7)? data_i[28] : 
                      (N9)? data_i[92] : 
                      (N11)? data_i[156] : 
                      (N13)? data_i[220] : 
                      (N8)? data_i[284] : 
                      (N10)? data_i[348] : 
                      (N12)? data_i[412] : 
                      (N14)? data_i[476] : 1'b0;
  assign data_o[27] = (N7)? data_i[27] : 
                      (N9)? data_i[91] : 
                      (N11)? data_i[155] : 
                      (N13)? data_i[219] : 
                      (N8)? data_i[283] : 
                      (N10)? data_i[347] : 
                      (N12)? data_i[411] : 
                      (N14)? data_i[475] : 1'b0;
  assign data_o[26] = (N7)? data_i[26] : 
                      (N9)? data_i[90] : 
                      (N11)? data_i[154] : 
                      (N13)? data_i[218] : 
                      (N8)? data_i[282] : 
                      (N10)? data_i[346] : 
                      (N12)? data_i[410] : 
                      (N14)? data_i[474] : 1'b0;
  assign data_o[25] = (N7)? data_i[25] : 
                      (N9)? data_i[89] : 
                      (N11)? data_i[153] : 
                      (N13)? data_i[217] : 
                      (N8)? data_i[281] : 
                      (N10)? data_i[345] : 
                      (N12)? data_i[409] : 
                      (N14)? data_i[473] : 1'b0;
  assign data_o[24] = (N7)? data_i[24] : 
                      (N9)? data_i[88] : 
                      (N11)? data_i[152] : 
                      (N13)? data_i[216] : 
                      (N8)? data_i[280] : 
                      (N10)? data_i[344] : 
                      (N12)? data_i[408] : 
                      (N14)? data_i[472] : 1'b0;
  assign data_o[23] = (N7)? data_i[23] : 
                      (N9)? data_i[87] : 
                      (N11)? data_i[151] : 
                      (N13)? data_i[215] : 
                      (N8)? data_i[279] : 
                      (N10)? data_i[343] : 
                      (N12)? data_i[407] : 
                      (N14)? data_i[471] : 1'b0;
  assign data_o[22] = (N7)? data_i[22] : 
                      (N9)? data_i[86] : 
                      (N11)? data_i[150] : 
                      (N13)? data_i[214] : 
                      (N8)? data_i[278] : 
                      (N10)? data_i[342] : 
                      (N12)? data_i[406] : 
                      (N14)? data_i[470] : 1'b0;
  assign data_o[21] = (N7)? data_i[21] : 
                      (N9)? data_i[85] : 
                      (N11)? data_i[149] : 
                      (N13)? data_i[213] : 
                      (N8)? data_i[277] : 
                      (N10)? data_i[341] : 
                      (N12)? data_i[405] : 
                      (N14)? data_i[469] : 1'b0;
  assign data_o[20] = (N7)? data_i[20] : 
                      (N9)? data_i[84] : 
                      (N11)? data_i[148] : 
                      (N13)? data_i[212] : 
                      (N8)? data_i[276] : 
                      (N10)? data_i[340] : 
                      (N12)? data_i[404] : 
                      (N14)? data_i[468] : 1'b0;
  assign data_o[19] = (N7)? data_i[19] : 
                      (N9)? data_i[83] : 
                      (N11)? data_i[147] : 
                      (N13)? data_i[211] : 
                      (N8)? data_i[275] : 
                      (N10)? data_i[339] : 
                      (N12)? data_i[403] : 
                      (N14)? data_i[467] : 1'b0;
  assign data_o[18] = (N7)? data_i[18] : 
                      (N9)? data_i[82] : 
                      (N11)? data_i[146] : 
                      (N13)? data_i[210] : 
                      (N8)? data_i[274] : 
                      (N10)? data_i[338] : 
                      (N12)? data_i[402] : 
                      (N14)? data_i[466] : 1'b0;
  assign data_o[17] = (N7)? data_i[17] : 
                      (N9)? data_i[81] : 
                      (N11)? data_i[145] : 
                      (N13)? data_i[209] : 
                      (N8)? data_i[273] : 
                      (N10)? data_i[337] : 
                      (N12)? data_i[401] : 
                      (N14)? data_i[465] : 1'b0;
  assign data_o[16] = (N7)? data_i[16] : 
                      (N9)? data_i[80] : 
                      (N11)? data_i[144] : 
                      (N13)? data_i[208] : 
                      (N8)? data_i[272] : 
                      (N10)? data_i[336] : 
                      (N12)? data_i[400] : 
                      (N14)? data_i[464] : 1'b0;
  assign data_o[15] = (N7)? data_i[15] : 
                      (N9)? data_i[79] : 
                      (N11)? data_i[143] : 
                      (N13)? data_i[207] : 
                      (N8)? data_i[271] : 
                      (N10)? data_i[335] : 
                      (N12)? data_i[399] : 
                      (N14)? data_i[463] : 1'b0;
  assign data_o[14] = (N7)? data_i[14] : 
                      (N9)? data_i[78] : 
                      (N11)? data_i[142] : 
                      (N13)? data_i[206] : 
                      (N8)? data_i[270] : 
                      (N10)? data_i[334] : 
                      (N12)? data_i[398] : 
                      (N14)? data_i[462] : 1'b0;
  assign data_o[13] = (N7)? data_i[13] : 
                      (N9)? data_i[77] : 
                      (N11)? data_i[141] : 
                      (N13)? data_i[205] : 
                      (N8)? data_i[269] : 
                      (N10)? data_i[333] : 
                      (N12)? data_i[397] : 
                      (N14)? data_i[461] : 1'b0;
  assign data_o[12] = (N7)? data_i[12] : 
                      (N9)? data_i[76] : 
                      (N11)? data_i[140] : 
                      (N13)? data_i[204] : 
                      (N8)? data_i[268] : 
                      (N10)? data_i[332] : 
                      (N12)? data_i[396] : 
                      (N14)? data_i[460] : 1'b0;
  assign data_o[11] = (N7)? data_i[11] : 
                      (N9)? data_i[75] : 
                      (N11)? data_i[139] : 
                      (N13)? data_i[203] : 
                      (N8)? data_i[267] : 
                      (N10)? data_i[331] : 
                      (N12)? data_i[395] : 
                      (N14)? data_i[459] : 1'b0;
  assign data_o[10] = (N7)? data_i[10] : 
                      (N9)? data_i[74] : 
                      (N11)? data_i[138] : 
                      (N13)? data_i[202] : 
                      (N8)? data_i[266] : 
                      (N10)? data_i[330] : 
                      (N12)? data_i[394] : 
                      (N14)? data_i[458] : 1'b0;
  assign data_o[9] = (N7)? data_i[9] : 
                     (N9)? data_i[73] : 
                     (N11)? data_i[137] : 
                     (N13)? data_i[201] : 
                     (N8)? data_i[265] : 
                     (N10)? data_i[329] : 
                     (N12)? data_i[393] : 
                     (N14)? data_i[457] : 1'b0;
  assign data_o[8] = (N7)? data_i[8] : 
                     (N9)? data_i[72] : 
                     (N11)? data_i[136] : 
                     (N13)? data_i[200] : 
                     (N8)? data_i[264] : 
                     (N10)? data_i[328] : 
                     (N12)? data_i[392] : 
                     (N14)? data_i[456] : 1'b0;
  assign data_o[7] = (N7)? data_i[7] : 
                     (N9)? data_i[71] : 
                     (N11)? data_i[135] : 
                     (N13)? data_i[199] : 
                     (N8)? data_i[263] : 
                     (N10)? data_i[327] : 
                     (N12)? data_i[391] : 
                     (N14)? data_i[455] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] : 
                     (N9)? data_i[70] : 
                     (N11)? data_i[134] : 
                     (N13)? data_i[198] : 
                     (N8)? data_i[262] : 
                     (N10)? data_i[326] : 
                     (N12)? data_i[390] : 
                     (N14)? data_i[454] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] : 
                     (N9)? data_i[69] : 
                     (N11)? data_i[133] : 
                     (N13)? data_i[197] : 
                     (N8)? data_i[261] : 
                     (N10)? data_i[325] : 
                     (N12)? data_i[389] : 
                     (N14)? data_i[453] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] : 
                     (N9)? data_i[68] : 
                     (N11)? data_i[132] : 
                     (N13)? data_i[196] : 
                     (N8)? data_i[260] : 
                     (N10)? data_i[324] : 
                     (N12)? data_i[388] : 
                     (N14)? data_i[452] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] : 
                     (N9)? data_i[67] : 
                     (N11)? data_i[131] : 
                     (N13)? data_i[195] : 
                     (N8)? data_i[259] : 
                     (N10)? data_i[323] : 
                     (N12)? data_i[387] : 
                     (N14)? data_i[451] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] : 
                     (N9)? data_i[66] : 
                     (N11)? data_i[130] : 
                     (N13)? data_i[194] : 
                     (N8)? data_i[258] : 
                     (N10)? data_i[322] : 
                     (N12)? data_i[386] : 
                     (N14)? data_i[450] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] : 
                     (N9)? data_i[65] : 
                     (N11)? data_i[129] : 
                     (N13)? data_i[193] : 
                     (N8)? data_i[257] : 
                     (N10)? data_i[321] : 
                     (N12)? data_i[385] : 
                     (N14)? data_i[449] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] : 
                     (N9)? data_i[64] : 
                     (N11)? data_i[128] : 
                     (N13)? data_i[192] : 
                     (N8)? data_i[256] : 
                     (N10)? data_i[320] : 
                     (N12)? data_i[384] : 
                     (N14)? data_i[448] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];

endmodule



module bsg_mux_width_p32_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [0:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[63] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[62] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[61] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[60] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[59] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[58] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[57] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[56] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[55] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[54] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[53] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[52] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[51] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[50] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[49] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[48] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[47] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[46] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[45] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[44] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[43] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[42] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[41] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[40] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[39] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[38] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[37] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[36] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[35] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[34] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[33] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[32] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_width_p16_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [1:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N4)? data_i[31] : 
                      (N3)? data_i[47] : 
                      (N5)? data_i[63] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N4)? data_i[30] : 
                      (N3)? data_i[46] : 
                      (N5)? data_i[62] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N4)? data_i[29] : 
                      (N3)? data_i[45] : 
                      (N5)? data_i[61] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N4)? data_i[28] : 
                      (N3)? data_i[44] : 
                      (N5)? data_i[60] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N4)? data_i[27] : 
                      (N3)? data_i[43] : 
                      (N5)? data_i[59] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N4)? data_i[26] : 
                      (N3)? data_i[42] : 
                      (N5)? data_i[58] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N4)? data_i[25] : 
                     (N3)? data_i[41] : 
                     (N5)? data_i[57] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N4)? data_i[24] : 
                     (N3)? data_i[40] : 
                     (N5)? data_i[56] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[23] : 
                     (N3)? data_i[39] : 
                     (N5)? data_i[55] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[22] : 
                     (N3)? data_i[38] : 
                     (N5)? data_i[54] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[21] : 
                     (N3)? data_i[37] : 
                     (N5)? data_i[53] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[20] : 
                     (N3)? data_i[36] : 
                     (N5)? data_i[52] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[19] : 
                     (N3)? data_i[35] : 
                     (N5)? data_i[51] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[18] : 
                     (N3)? data_i[34] : 
                     (N5)? data_i[50] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[17] : 
                     (N3)? data_i[33] : 
                     (N5)? data_i[49] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[16] : 
                     (N3)? data_i[32] : 
                     (N5)? data_i[48] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p8_els_p8
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [2:0] sel_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  assign data_o[7] = (N7)? data_i[7] : 
                     (N9)? data_i[15] : 
                     (N11)? data_i[23] : 
                     (N13)? data_i[31] : 
                     (N8)? data_i[39] : 
                     (N10)? data_i[47] : 
                     (N12)? data_i[55] : 
                     (N14)? data_i[63] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] : 
                     (N9)? data_i[14] : 
                     (N11)? data_i[22] : 
                     (N13)? data_i[30] : 
                     (N8)? data_i[38] : 
                     (N10)? data_i[46] : 
                     (N12)? data_i[54] : 
                     (N14)? data_i[62] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] : 
                     (N9)? data_i[13] : 
                     (N11)? data_i[21] : 
                     (N13)? data_i[29] : 
                     (N8)? data_i[37] : 
                     (N10)? data_i[45] : 
                     (N12)? data_i[53] : 
                     (N14)? data_i[61] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] : 
                     (N9)? data_i[12] : 
                     (N11)? data_i[20] : 
                     (N13)? data_i[28] : 
                     (N8)? data_i[36] : 
                     (N10)? data_i[44] : 
                     (N12)? data_i[52] : 
                     (N14)? data_i[60] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] : 
                     (N9)? data_i[11] : 
                     (N11)? data_i[19] : 
                     (N13)? data_i[27] : 
                     (N8)? data_i[35] : 
                     (N10)? data_i[43] : 
                     (N12)? data_i[51] : 
                     (N14)? data_i[59] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] : 
                     (N9)? data_i[10] : 
                     (N11)? data_i[18] : 
                     (N13)? data_i[26] : 
                     (N8)? data_i[34] : 
                     (N10)? data_i[42] : 
                     (N12)? data_i[50] : 
                     (N14)? data_i[58] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] : 
                     (N9)? data_i[9] : 
                     (N11)? data_i[17] : 
                     (N13)? data_i[25] : 
                     (N8)? data_i[33] : 
                     (N10)? data_i[41] : 
                     (N12)? data_i[49] : 
                     (N14)? data_i[57] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] : 
                     (N9)? data_i[8] : 
                     (N11)? data_i[16] : 
                     (N13)? data_i[24] : 
                     (N8)? data_i[32] : 
                     (N10)? data_i[40] : 
                     (N12)? data_i[48] : 
                     (N14)? data_i[56] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];

endmodule



module bsg_decode_num_out_p8
(
  i,
  o
);

  input [2:0] i;
  output [7:0] o;
  wire [7:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bp_be_dcache_lru_decode_ways_p8
(
  way_id_i,
  data_o,
  mask_o
);

  input [2:0] way_id_i;
  output [6:0] data_o;
  output [6:0] mask_o;
  wire [6:0] data_o,mask_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30;
  assign mask_o[0] = 1'b1;
  assign N11 = N8 & N9;
  assign N12 = N11 & N10;
  assign N13 = way_id_i[2] | way_id_i[1];
  assign N14 = N13 | N10;
  assign N16 = way_id_i[2] | N9;
  assign N17 = N16 | way_id_i[0];
  assign N19 = N16 | N10;
  assign N21 = N8 | way_id_i[1];
  assign N22 = N21 | way_id_i[0];
  assign N24 = N21 | N10;
  assign N26 = N8 | N9;
  assign N27 = N26 | way_id_i[0];
  assign N29 = way_id_i[2] & way_id_i[1];
  assign N30 = N29 & way_id_i[0];
  assign data_o = (N0)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                  (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                  (N2)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                  (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                  (N4)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                  (N6)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                  (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N12;
  assign N1 = N15;
  assign N2 = N18;
  assign N3 = N20;
  assign N4 = N23;
  assign N5 = N25;
  assign N6 = N28;
  assign N7 = N30;
  assign mask_o[6:1] = (N0)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                       (N1)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                       (N2)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                       (N3)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                       (N4)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                       (N5)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                       (N6)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                       (N7)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 1'b0;
  assign N8 = ~way_id_i[2];
  assign N9 = ~way_id_i[1];
  assign N10 = ~way_id_i[0];
  assign N15 = ~N14;
  assign N18 = ~N17;
  assign N20 = ~N19;
  assign N23 = ~N22;
  assign N25 = ~N24;
  assign N28 = ~N27;

endmodule



module bsg_decode_with_v_num_out_p8
(
  i,
  v_i,
  o
);

  input [2:0] i;
  output [7:0] o;
  input v_i;
  wire [7:0] o,lo;

  bsg_decode_num_out_p8
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bp_be_dcache_data_width_p64_paddr_width_p22_sets_p64_ways_p8_num_cce_p1_num_lce_p2
(
  clk_i,
  reset_i,
  lce_id_i,
  dcache_pkt_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  tlb_miss_i,
  ptag_i,
  cache_miss_o,
  poison_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_tr_resp_i,
  lce_tr_resp_v_i,
  lce_tr_resp_ready_o,
  lce_tr_resp_o,
  lce_tr_resp_v_o,
  lce_tr_resp_ready_i
);

  input [0:0] lce_id_i;
  input [79:0] dcache_pkt_i;
  output [63:0] data_o;
  input [9:0] ptag_i;
  output [29:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [539:0] lce_data_cmd_i;
  input [538:0] lce_tr_resp_i;
  output [538:0] lce_tr_resp_o;
  input clk_i;
  input reset_i;
  input v_i;
  input tlb_miss_i;
  input poison_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_tr_resp_v_i;
  input lce_tr_resp_ready_i;
  output ready_o;
  output v_o;
  output cache_miss_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_tr_resp_ready_o;
  output lce_tr_resp_v_o;
  wire [63:0] data_o,data_mem_mask_li,bypass_data_lo,ld_data_way_picked,bypass_data_masked;
  wire [29:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [538:0] lce_tr_resp_o;
  wire ready_o,v_o,cache_miss_o,lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,
  lce_cmd_ready_o,lce_data_cmd_ready_o,lce_tr_resp_ready_o,lce_tr_resp_v_o,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,load_op,
  signed_op,tl_we,N65,N66,N67,N68,N69,N70,n_0_net_,tag_mem_w_li,tag_mem_v_li,
  n_1_net_,n_2_net_,n_3_net_,n_4_net_,n_5_net_,n_6_net_,n_7_net_,n_8_net_,tv_we,N71,N72,
  N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,N100,load_hit,store_hit,load_miss_tv,store_miss_tv,
  wbuf_v_li,wbuf_entry_in_data__63_,wbuf_entry_in_data__62_,
  wbuf_entry_in_data__61_,wbuf_entry_in_data__60_,wbuf_entry_in_data__59_,wbuf_entry_in_data__58_,
  wbuf_entry_in_data__57_,wbuf_entry_in_data__56_,wbuf_entry_in_data__55_,
  wbuf_entry_in_data__54_,wbuf_entry_in_data__53_,wbuf_entry_in_data__52_,
  wbuf_entry_in_data__51_,wbuf_entry_in_data__50_,wbuf_entry_in_data__49_,wbuf_entry_in_data__48_,
  wbuf_entry_in_data__47_,wbuf_entry_in_data__46_,wbuf_entry_in_data__45_,
  wbuf_entry_in_data__44_,wbuf_entry_in_data__43_,wbuf_entry_in_data__42_,
  wbuf_entry_in_data__41_,wbuf_entry_in_data__40_,wbuf_entry_in_data__39_,wbuf_entry_in_data__38_,
  wbuf_entry_in_data__37_,wbuf_entry_in_data__36_,wbuf_entry_in_data__35_,
  wbuf_entry_in_data__34_,wbuf_entry_in_data__33_,wbuf_entry_in_data__32_,
  wbuf_entry_in_data__31_,wbuf_entry_in_data__30_,wbuf_entry_in_data__29_,wbuf_entry_in_data__28_,
  wbuf_entry_in_data__27_,wbuf_entry_in_data__26_,wbuf_entry_in_data__25_,
  wbuf_entry_in_data__24_,wbuf_entry_in_data__23_,wbuf_entry_in_data__22_,
  wbuf_entry_in_data__21_,wbuf_entry_in_data__20_,wbuf_entry_in_data__19_,wbuf_entry_in_data__18_,
  wbuf_entry_in_data__17_,wbuf_entry_in_data__16_,wbuf_entry_in_data__15_,
  wbuf_entry_in_data__14_,wbuf_entry_in_data__13_,wbuf_entry_in_data__12_,
  wbuf_entry_in_data__11_,wbuf_entry_in_data__10_,wbuf_entry_in_data__9_,wbuf_entry_in_data__8_,
  wbuf_entry_in_mask__7_,wbuf_entry_in_mask__6_,wbuf_entry_in_mask__5_,
  wbuf_entry_in_mask__4_,wbuf_entry_in_mask__3_,wbuf_entry_in_mask__2_,wbuf_entry_in_mask__1_,
  wbuf_entry_in_mask__0_,wbuf_v_lo,wbuf_yumi_li,wbuf_empty_lo,bypass_v_li,
  lce_snoop_match_lo,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,n_10_net_,stat_mem_w_li,stat_mem_v_li,invalid_exist,N135,
  lce_data_mem_pkt_v_lo,lce_data_mem_pkt_yumi_li,lce_tag_mem_pkt_v_lo,
  lce_tag_mem_pkt_yumi_li,lce_stat_mem_pkt_v_lo,lce_stat_mem_pkt_yumi_li,n_13_net__2_,n_13_net__1_,
  n_13_net__0_,genblk4_word_sigext,genblk4_half_sigext,genblk4_byte_sigext,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,n_14_net__2_,n_14_net__1_,n_14_net__0_,N207,N208,N209,
  N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,
  N226,N227,N228,N229,n_18_net__0_,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,
  N240,n_20_net__1_,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,
  n_22_net__1_,n_22_net__0_,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,
  n_24_net__2_,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  n_26_net__2_,n_26_net__0_,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,
  n_28_net__2_,n_28_net__1_,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,
  N299,N300,n_30_net__2_,n_30_net__1_,n_30_net__0_,N301,N302,N303,N304,N305,N306,
  N307,N308,N309,N310,N311,N312,N313,N314,N315,dirty_mask_v_li,N316,N317,N318,N319,
  N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,
  N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
  N352,N353,N354,N355,N356,n_33_net__0_,n_34_net__1_,n_35_net__1_,n_35_net__0_,
  n_36_net__2_,n_37_net__2_,n_37_net__0_,n_38_net__2_,n_38_net__1_,n_39_net__2_,
  n_39_net__1_,n_39_net__0_,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484;
  wire [5:0] tag_mem_addr_li,stat_mem_addr_li;
  wire [95:0] tag_mem_data_li,tag_mem_mask_li,tag_mem_data_lo;
  wire [7:0] data_mem_w_li,data_mem_v_li,load_hit_tv,store_hit_tv,bypass_mask_lo,
  genblk4_data_byte_selected,wbuf_data_mem_v,lce_tag_mem_way_one_hot,dirty_mask_lo;
  wire [71:0] data_mem_addr_li;
  wire [511:0] data_mem_data_li,data_mem_data_lo,lce_data_mem_data_li,lce_data_mem_write_data;
  wire [2:0] load_hit_way,store_hit_way,lru_encode,invalid_way,lce_lru_way_li,
  lru_decode_way_li,dirty_mask_way_li;
  wire [96:0] wbuf_entry_out;
  wire [14:0] stat_mem_data_li,stat_mem_mask_li,stat_mem_data_lo;
  wire [521:0] lce_data_mem_pkt;
  wire [22:0] lce_tag_mem_pkt;
  wire [10:0] lce_stat_mem_pkt;
  wire [31:0] genblk4_data_word_selected;
  wire [15:0] genblk4_data_half_selected;
  wire [6:0] lru_decode_data_lo,lru_decode_mask_lo;
  reg [63:0] data_tl_r,data_tv_r;
  reg v_tl_r,load_op_tl_r,store_op_tl_r,signed_op_tl_r,double_op_tl_r,word_op_tl_r,
  half_op_tl_r,v_tv_r,load_op_tv_r,store_op_tv_r,double_op_tv_r,signed_op_tv_r,
  word_op_tv_r,half_op_tv_r;
  reg [11:0] page_offset_tl_r;
  reg [95:0] tag_info_tv_r;
  reg [21:0] paddr_tv_r;
  reg [511:0] ld_data_tv_r;
  reg [2:0] lce_data_mem_pkt_way_r;

  bsg_mem_1rw_sync_mask_write_bit_width_p96_els_p64
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(n_0_net_),
    .w_mask_i(tag_mem_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_0__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_1_net_),
    .w_i(data_mem_w_li[0]),
    .addr_i(data_mem_addr_li[8:0]),
    .data_i(data_mem_data_li[63:0]),
    .write_mask_i(data_mem_mask_li[7:0]),
    .data_o(data_mem_data_lo[63:0])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_1__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_2_net_),
    .w_i(data_mem_w_li[1]),
    .addr_i(data_mem_addr_li[17:9]),
    .data_i(data_mem_data_li[127:64]),
    .write_mask_i(data_mem_mask_li[15:8]),
    .data_o(data_mem_data_lo[127:64])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_2__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_3_net_),
    .w_i(data_mem_w_li[2]),
    .addr_i(data_mem_addr_li[26:18]),
    .data_i(data_mem_data_li[191:128]),
    .write_mask_i(data_mem_mask_li[23:16]),
    .data_o(data_mem_data_lo[191:128])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_3__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_4_net_),
    .w_i(data_mem_w_li[3]),
    .addr_i(data_mem_addr_li[35:27]),
    .data_i(data_mem_data_li[255:192]),
    .write_mask_i(data_mem_mask_li[31:24]),
    .data_o(data_mem_data_lo[255:192])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_4__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_5_net_),
    .w_i(data_mem_w_li[4]),
    .addr_i(data_mem_addr_li[44:36]),
    .data_i(data_mem_data_li[319:256]),
    .write_mask_i(data_mem_mask_li[39:32]),
    .data_o(data_mem_data_lo[319:256])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_5__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_6_net_),
    .w_i(data_mem_w_li[5]),
    .addr_i(data_mem_addr_li[53:45]),
    .data_i(data_mem_data_li[383:320]),
    .write_mask_i(data_mem_mask_li[47:40]),
    .data_o(data_mem_data_lo[383:320])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_6__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_7_net_),
    .w_i(data_mem_w_li[6]),
    .addr_i(data_mem_addr_li[62:54]),
    .data_i(data_mem_data_li[447:384]),
    .write_mask_i(data_mem_mask_li[55:48]),
    .data_o(data_mem_data_lo[447:384])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_7__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_8_net_),
    .w_i(data_mem_w_li[7]),
    .addr_i(data_mem_addr_li[71:63]),
    .data_i(data_mem_data_li[511:448]),
    .write_mask_i(data_mem_mask_li[63:56]),
    .data_o(data_mem_data_lo[511:448])
  );

  assign N85 = paddr_tv_r[21:12] == tag_info_tv_r[9:0];
  assign N86 = paddr_tv_r[21:12] == tag_info_tv_r[9:0];
  assign N87 = paddr_tv_r[21:12] == tag_info_tv_r[21:12];
  assign N88 = paddr_tv_r[21:12] == tag_info_tv_r[21:12];
  assign N89 = paddr_tv_r[21:12] == tag_info_tv_r[33:24];
  assign N90 = paddr_tv_r[21:12] == tag_info_tv_r[33:24];
  assign N91 = paddr_tv_r[21:12] == tag_info_tv_r[45:36];
  assign N92 = paddr_tv_r[21:12] == tag_info_tv_r[45:36];
  assign N93 = paddr_tv_r[21:12] == tag_info_tv_r[57:48];
  assign N94 = paddr_tv_r[21:12] == tag_info_tv_r[57:48];
  assign N95 = paddr_tv_r[21:12] == tag_info_tv_r[69:60];
  assign N96 = paddr_tv_r[21:12] == tag_info_tv_r[69:60];
  assign N97 = paddr_tv_r[21:12] == tag_info_tv_r[81:72];
  assign N98 = paddr_tv_r[21:12] == tag_info_tv_r[81:72];
  assign N99 = paddr_tv_r[21:12] == tag_info_tv_r[93:84];
  assign N100 = paddr_tv_r[21:12] == tag_info_tv_r[93:84];

  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_load_hit
  (
    .i(load_hit_tv),
    .addr_o(load_hit_way),
    .v_o(load_hit)
  );


  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_store_hit
  (
    .i(store_hit_tv),
    .addr_o(store_hit_way),
    .v_o(store_hit)
  );


  bp_be_dcache_wbuf_data_width_p64_paddr_width_p22_ways_p8_sets_p64
  wbuf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(wbuf_v_li),
    .wbuf_entry_i({ paddr_tv_r, wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_, data_tv_r[7:0], wbuf_entry_in_mask__7_, wbuf_entry_in_mask__6_, wbuf_entry_in_mask__5_, wbuf_entry_in_mask__4_, wbuf_entry_in_mask__3_, wbuf_entry_in_mask__2_, wbuf_entry_in_mask__1_, wbuf_entry_in_mask__0_, store_hit_way }),
    .yumi_i(wbuf_yumi_li),
    .v_o(wbuf_v_lo),
    .wbuf_entry_o(wbuf_entry_out),
    .empty_o(wbuf_empty_lo),
    .bypass_addr_i({ ptag_i, page_offset_tl_r }),
    .bypass_v_i(bypass_v_li),
    .bypass_data_o(bypass_data_lo),
    .bypass_mask_o(bypass_mask_lo),
    .lce_snoop_index_i(lce_data_mem_pkt[521:516]),
    .lce_snoop_way_i(lce_data_mem_pkt[515:513]),
    .lce_snoop_match_o(lce_snoop_match_lo)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p15_els_p64
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(n_10_net_),
    .w_mask_i(stat_mem_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_data_lo)
  );


  bp_be_dcache_lru_encode_ways_p8
  lru_encoder
  (
    .lru_i(stat_mem_data_lo[14:8]),
    .way_id_o(lru_encode)
  );


  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_invalid
  (
    .i({ N358, N360, N362, N364, N366, N368, N370, N372 }),
    .addr_o(invalid_way),
    .v_o(invalid_exist)
  );


  bp_be_dcache_lce_data_width_p64_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_num_cce_p1_num_lce_p2
  lce
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_id_i(lce_id_i[0]),
    .ready_o(ready_o),
    .cache_miss_o(cache_miss_o),
    .load_miss_i(load_miss_tv),
    .store_miss_i(store_miss_tv),
    .miss_addr_i(paddr_tv_r),
    .data_mem_pkt_v_o(lce_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_data_mem_pkt),
    .data_mem_data_i(lce_data_mem_data_li),
    .data_mem_pkt_yumi_i(lce_data_mem_pkt_yumi_li),
    .tag_mem_pkt_v_o(lce_tag_mem_pkt_v_lo),
    .tag_mem_pkt_o(lce_tag_mem_pkt),
    .tag_mem_pkt_yumi_i(lce_tag_mem_pkt_yumi_li),
    .stat_mem_pkt_v_o(lce_stat_mem_pkt_v_lo),
    .stat_mem_pkt_o(lce_stat_mem_pkt),
    .lru_way_i(lce_lru_way_li),
    .dirty_i(stat_mem_data_lo[7:0]),
    .stat_mem_pkt_yumi_i(lce_stat_mem_pkt_yumi_li),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_tr_resp_i(lce_tr_resp_i),
    .lce_tr_resp_v_i(lce_tr_resp_v_i),
    .lce_tr_resp_ready_o(lce_tr_resp_ready_o),
    .lce_tr_resp_o(lce_tr_resp_o),
    .lce_tr_resp_v_o(lce_tr_resp_v_o),
    .lce_tr_resp_ready_i(lce_tr_resp_ready_i)
  );


  bsg_mux_width_p64_els_p8
  ld_data_set_select_mux
  (
    .data_i(ld_data_tv_r),
    .sel_i({ n_13_net__2_, n_13_net__1_, n_13_net__0_ }),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_segmented_segments_p8_segment_width_p8
  bypass_mux_segmented
  (
    .data0_i(ld_data_way_picked),
    .data1_i(bypass_data_lo),
    .sel_i(bypass_mask_lo),
    .data_o(bypass_data_masked)
  );


  bsg_mux_width_p32_els_p2
  genblk4_word_mux
  (
    .data_i(bypass_data_masked),
    .sel_i(paddr_tv_r[2]),
    .data_o(genblk4_data_word_selected)
  );


  bsg_mux_width_p16_els_p4
  genblk4_half_mux
  (
    .data_i(bypass_data_masked),
    .sel_i(paddr_tv_r[2:1]),
    .data_o(genblk4_data_half_selected)
  );


  bsg_mux_width_p8_els_p8
  genblk4_byte_mux
  (
    .data_i(bypass_data_masked),
    .sel_i(paddr_tv_r[2:0]),
    .data_o(genblk4_data_byte_selected)
  );


  bsg_decode_num_out_p8
  wbuf_data_mem_v_decode
  (
    .i({ n_14_net__2_, n_14_net__1_, n_14_net__0_ }),
    .o(wbuf_data_mem_v)
  );


  bsg_mux_width_p64_els_p8
  genblk5_0__lce_data_mem_write_mux
  (
    .data_i(lce_data_mem_pkt[512:1]),
    .sel_i(lce_data_mem_pkt[515:513]),
    .data_o(lce_data_mem_write_data[63:0])
  );


  bsg_mux_width_p64_els_p8
  genblk5_1__lce_data_mem_write_mux
  (
    .data_i(lce_data_mem_pkt[512:1]),
    .sel_i({ lce_data_mem_pkt[515:514], n_18_net__0_ }),
    .data_o(lce_data_mem_write_data[127:64])
  );


  bsg_mux_width_p64_els_p8
  genblk5_2__lce_data_mem_write_mux
  (
    .data_i(lce_data_mem_pkt[512:1]),
    .sel_i({ lce_data_mem_pkt[515:515], n_20_net__1_, lce_data_mem_pkt[513:513] }),
    .data_o(lce_data_mem_write_data[191:128])
  );


  bsg_mux_width_p64_els_p8
  genblk5_3__lce_data_mem_write_mux
  (
    .data_i(lce_data_mem_pkt[512:1]),
    .sel_i({ lce_data_mem_pkt[515:515], n_22_net__1_, n_22_net__0_ }),
    .data_o(lce_data_mem_write_data[255:192])
  );


  bsg_mux_width_p64_els_p8
  genblk5_4__lce_data_mem_write_mux
  (
    .data_i(lce_data_mem_pkt[512:1]),
    .sel_i({ n_24_net__2_, lce_data_mem_pkt[514:513] }),
    .data_o(lce_data_mem_write_data[319:256])
  );


  bsg_mux_width_p64_els_p8
  genblk5_5__lce_data_mem_write_mux
  (
    .data_i(lce_data_mem_pkt[512:1]),
    .sel_i({ n_26_net__2_, lce_data_mem_pkt[514:514], n_26_net__0_ }),
    .data_o(lce_data_mem_write_data[383:320])
  );


  bsg_mux_width_p64_els_p8
  genblk5_6__lce_data_mem_write_mux
  (
    .data_i(lce_data_mem_pkt[512:1]),
    .sel_i({ n_28_net__2_, n_28_net__1_, lce_data_mem_pkt[513:513] }),
    .data_o(lce_data_mem_write_data[447:384])
  );


  bsg_mux_width_p64_els_p8
  genblk5_7__lce_data_mem_write_mux
  (
    .data_i(lce_data_mem_pkt[512:1]),
    .sel_i({ n_30_net__2_, n_30_net__1_, n_30_net__0_ }),
    .data_o(lce_data_mem_write_data[511:448])
  );


  bsg_decode_num_out_p8
  lce_tag_mem_way_decode
  (
    .i(lce_tag_mem_pkt[16:14]),
    .o(lce_tag_mem_way_one_hot)
  );

  assign N307 = N305 & N306;
  assign N308 = lce_tag_mem_pkt[1] | N306;
  assign N310 = N305 | lce_tag_mem_pkt[0];
  assign N312 = lce_tag_mem_pkt[1] & lce_tag_mem_pkt[0];

  bp_be_dcache_lru_decode_ways_p8
  lru_decode
  (
    .way_id_i(lru_decode_way_li),
    .data_o(lru_decode_data_lo),
    .mask_o(lru_decode_mask_lo)
  );


  bsg_decode_with_v_num_out_p8
  dirty_mask_decode
  (
    .i(dirty_mask_way_li),
    .v_i(dirty_mask_v_li),
    .o(dirty_mask_lo)
  );

  assign N321 = N320 & N405;
  assign N322 = N320 | lce_stat_mem_pkt[0];
  assign N324 = lce_stat_mem_pkt[1] & lce_stat_mem_pkt[0];
  assign N325 = lce_stat_mem_pkt[1] | N405;

  bsg_mux_width_p64_els_p8
  genblk6_0__lce_data_mem_read_mux
  (
    .data_i(data_mem_data_lo),
    .sel_i(lce_data_mem_pkt_way_r),
    .data_o(lce_data_mem_data_li[63:0])
  );


  bsg_mux_width_p64_els_p8
  genblk6_1__lce_data_mem_read_mux
  (
    .data_i(data_mem_data_lo),
    .sel_i({ lce_data_mem_pkt_way_r[2:1], n_33_net__0_ }),
    .data_o(lce_data_mem_data_li[127:64])
  );


  bsg_mux_width_p64_els_p8
  genblk6_2__lce_data_mem_read_mux
  (
    .data_i(data_mem_data_lo),
    .sel_i({ lce_data_mem_pkt_way_r[2:2], n_34_net__1_, lce_data_mem_pkt_way_r[0:0] }),
    .data_o(lce_data_mem_data_li[191:128])
  );


  bsg_mux_width_p64_els_p8
  genblk6_3__lce_data_mem_read_mux
  (
    .data_i(data_mem_data_lo),
    .sel_i({ lce_data_mem_pkt_way_r[2:2], n_35_net__1_, n_35_net__0_ }),
    .data_o(lce_data_mem_data_li[255:192])
  );


  bsg_mux_width_p64_els_p8
  genblk6_4__lce_data_mem_read_mux
  (
    .data_i(data_mem_data_lo),
    .sel_i({ n_36_net__2_, lce_data_mem_pkt_way_r[1:0] }),
    .data_o(lce_data_mem_data_li[319:256])
  );


  bsg_mux_width_p64_els_p8
  genblk6_5__lce_data_mem_read_mux
  (
    .data_i(data_mem_data_lo),
    .sel_i({ n_37_net__2_, lce_data_mem_pkt_way_r[1:1], n_37_net__0_ }),
    .data_o(lce_data_mem_data_li[383:320])
  );


  bsg_mux_width_p64_els_p8
  genblk6_6__lce_data_mem_read_mux
  (
    .data_i(data_mem_data_lo),
    .sel_i({ n_38_net__2_, n_38_net__1_, lce_data_mem_pkt_way_r[0:0] }),
    .data_o(lce_data_mem_data_li[447:384])
  );


  bsg_mux_width_p64_els_p8
  genblk6_7__lce_data_mem_read_mux
  (
    .data_i(data_mem_data_lo),
    .sel_i({ n_39_net__2_, n_39_net__1_, n_39_net__0_ }),
    .data_o(lce_data_mem_data_li[511:448])
  );

  assign N357 = tag_info_tv_r[94] | tag_info_tv_r[95];
  assign N358 = ~N357;
  assign N359 = tag_info_tv_r[82] | tag_info_tv_r[83];
  assign N360 = ~N359;
  assign N361 = tag_info_tv_r[70] | tag_info_tv_r[71];
  assign N362 = ~N361;
  assign N363 = tag_info_tv_r[58] | tag_info_tv_r[59];
  assign N364 = ~N363;
  assign N365 = tag_info_tv_r[46] | tag_info_tv_r[47];
  assign N366 = ~N365;
  assign N367 = tag_info_tv_r[34] | tag_info_tv_r[35];
  assign N368 = ~N367;
  assign N369 = tag_info_tv_r[22] | tag_info_tv_r[23];
  assign N370 = ~N369;
  assign N371 = tag_info_tv_r[10] | tag_info_tv_r[11];
  assign N372 = ~N371;
  assign N373 = tag_info_tv_r[94] | tag_info_tv_r[95];
  assign N374 = tag_info_tv_r[82] | tag_info_tv_r[83];
  assign N375 = tag_info_tv_r[70] | tag_info_tv_r[71];
  assign N376 = tag_info_tv_r[58] | tag_info_tv_r[59];
  assign N377 = tag_info_tv_r[46] | tag_info_tv_r[47];
  assign N378 = tag_info_tv_r[34] | tag_info_tv_r[35];
  assign N379 = tag_info_tv_r[22] | tag_info_tv_r[23];
  assign N380 = tag_info_tv_r[10] | tag_info_tv_r[11];
  assign N381 = ~tag_info_tv_r[95];
  assign N382 = tag_info_tv_r[94] | N381;
  assign N383 = ~N382;
  assign N384 = ~tag_info_tv_r[83];
  assign N385 = tag_info_tv_r[82] | N384;
  assign N386 = ~N385;
  assign N387 = ~tag_info_tv_r[71];
  assign N388 = tag_info_tv_r[70] | N387;
  assign N389 = ~N388;
  assign N390 = ~tag_info_tv_r[59];
  assign N391 = tag_info_tv_r[58] | N390;
  assign N392 = ~N391;
  assign N393 = ~tag_info_tv_r[47];
  assign N394 = tag_info_tv_r[46] | N393;
  assign N395 = ~N394;
  assign N396 = ~tag_info_tv_r[35];
  assign N397 = tag_info_tv_r[34] | N396;
  assign N398 = ~N397;
  assign N399 = ~tag_info_tv_r[23];
  assign N400 = tag_info_tv_r[22] | N399;
  assign N401 = ~N400;
  assign N402 = ~tag_info_tv_r[11];
  assign N403 = tag_info_tv_r[10] | N402;
  assign N404 = ~N403;
  assign N405 = ~lce_stat_mem_pkt[0];
  assign N406 = N405 | lce_stat_mem_pkt[1];
  assign N407 = dcache_pkt_i[76] & dcache_pkt_i[77];
  assign N408 = ~dcache_pkt_i[77];
  assign N409 = dcache_pkt_i[76] | N408;
  assign N410 = ~N409;
  assign N411 = ~dcache_pkt_i[76];
  assign N412 = N411 | dcache_pkt_i[77];
  assign N413 = ~N412;
  assign N68 = (N0)? 1'b0 : 
               (N1)? tl_we : 1'b0;
  assign N0 = N66;
  assign N1 = N65;
  assign N69 = (N0)? 1'b0 : 
               (N1)? tl_we : 1'b0;
  assign N70 = (N0)? 1'b0 : 
               (N1)? N67 : 1'b0;
  assign N75 = (N2)? 1'b0 : 
               (N3)? tv_we : 1'b0;
  assign N2 = N72;
  assign N3 = N71;
  assign N76 = (N2)? 1'b0 : 
               (N3)? tv_we : 1'b0;
  assign N77 = (N2)? 1'b0 : 
               (N3)? tv_we : 1'b0;
  assign { N83, N82, N81, N80, N79, N78 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N3)? { N73, N73, N73, N73, N73, N73 } : 1'b0;
  assign N84 = (N2)? 1'b0 : 
               (N3)? N74 : 1'b0;
  assign { wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_ } = (N4)? data_tv_r[63:8] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N105)? { data_tv_r[31:0], data_tv_r[31:8] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N108)? { data_tv_r[15:0], data_tv_r[15:0], data_tv_r[15:0], data_tv_r[15:8] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N103)? { data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0] } : 1'b0;
  assign N4 = double_op_tv_r;
  assign { wbuf_entry_in_mask__7_, wbuf_entry_in_mask__6_, wbuf_entry_in_mask__5_, wbuf_entry_in_mask__4_, wbuf_entry_in_mask__3_, wbuf_entry_in_mask__2_, wbuf_entry_in_mask__1_, wbuf_entry_in_mask__0_ } = (N4)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N132)? { paddr_tv_r[2:2], paddr_tv_r[2:2], paddr_tv_r[2:2], paddr_tv_r[2:2], N112, N113, N114, N115 } : 
                                                                                                                                                                                                              (N134)? { N116, N117, N118, N119, N120, N121, N122, N123 } : 
                                                                                                                                                                                                              (N111)? { N124, N125, N126, N127, N128, N129, N130, N131 } : 1'b0;
  assign lce_lru_way_li = (N5)? invalid_way : 
                          (N6)? lru_encode : 1'b0;
  assign N5 = invalid_exist;
  assign N6 = N135;
  assign { N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140 } = (N4)? bypass_data_masked : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N204)? { genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_data_word_selected } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N206)? { genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_data_half_selected } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N139)? { genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_data_byte_selected } : 1'b0;
  assign data_o = (N7)? { N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140 } : 
                  (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N7 = load_op_tv_r;
  assign N8 = N136;
  assign data_mem_v_li = (N9)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                         (N212)? wbuf_data_mem_v : 
                         (N210)? { lce_data_mem_pkt_yumi_li, lce_data_mem_pkt_yumi_li, lce_data_mem_pkt_yumi_li, lce_data_mem_pkt_yumi_li, lce_data_mem_pkt_yumi_li, lce_data_mem_pkt_yumi_li, lce_data_mem_pkt_yumi_li, lce_data_mem_pkt_yumi_li } : 1'b0;
  assign N9 = N207;
  assign data_mem_addr_li[8:0] = (N10)? dcache_pkt_i[75:67] : 
                                 (N218)? wbuf_entry_out[86:78] : 
                                 (N216)? lce_data_mem_pkt[521:513] : 1'b0;
  assign N10 = N213;
  assign data_mem_data_li[63:0] = (N11)? wbuf_entry_out[74:11] : 
                                  (N12)? lce_data_mem_write_data[63:0] : 1'b0;
  assign N11 = N220;
  assign N12 = N219;
  assign data_mem_mask_li[7:0] = (N13)? wbuf_entry_out[10:3] : 
                                 (N14)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N13 = N222;
  assign N14 = N221;
  assign data_mem_addr_li[17:9] = (N15)? dcache_pkt_i[75:67] : 
                                  (N229)? wbuf_entry_out[86:78] : 
                                  (N226)? { lce_data_mem_pkt[521:514], N227 } : 1'b0;
  assign N15 = N223;
  assign data_mem_data_li[127:64] = (N16)? wbuf_entry_out[74:11] : 
                                    (N17)? lce_data_mem_write_data[127:64] : 1'b0;
  assign N16 = N231;
  assign N17 = N230;
  assign data_mem_mask_li[15:8] = (N18)? wbuf_entry_out[10:3] : 
                                  (N19)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N18 = N233;
  assign N19 = N232;
  assign data_mem_addr_li[26:18] = (N20)? dcache_pkt_i[75:67] : 
                                   (N240)? wbuf_entry_out[86:78] : 
                                   (N237)? { lce_data_mem_pkt[521:515], N238, lce_data_mem_pkt[513:513] } : 1'b0;
  assign N20 = N234;
  assign data_mem_data_li[191:128] = (N21)? wbuf_entry_out[74:11] : 
                                     (N22)? lce_data_mem_write_data[191:128] : 1'b0;
  assign N21 = N242;
  assign N22 = N241;
  assign data_mem_mask_li[23:16] = (N23)? wbuf_entry_out[10:3] : 
                                   (N24)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N23 = N244;
  assign N24 = N243;
  assign data_mem_addr_li[35:27] = (N25)? dcache_pkt_i[75:67] : 
                                   (N252)? wbuf_entry_out[86:78] : 
                                   (N248)? { lce_data_mem_pkt[521:515], N249, N250 } : 1'b0;
  assign N25 = N245;
  assign data_mem_data_li[255:192] = (N26)? wbuf_entry_out[74:11] : 
                                     (N27)? lce_data_mem_write_data[255:192] : 1'b0;
  assign N26 = N254;
  assign N27 = N253;
  assign data_mem_mask_li[31:24] = (N28)? wbuf_entry_out[10:3] : 
                                   (N29)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N28 = N256;
  assign N29 = N255;
  assign data_mem_addr_li[44:36] = (N30)? dcache_pkt_i[75:67] : 
                                   (N263)? wbuf_entry_out[86:78] : 
                                   (N260)? { lce_data_mem_pkt[521:516], N261, lce_data_mem_pkt[514:513] } : 1'b0;
  assign N30 = N257;
  assign data_mem_data_li[319:256] = (N31)? wbuf_entry_out[74:11] : 
                                     (N32)? lce_data_mem_write_data[319:256] : 1'b0;
  assign N31 = N265;
  assign N32 = N264;
  assign data_mem_mask_li[39:32] = (N33)? wbuf_entry_out[10:3] : 
                                   (N34)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N33 = N267;
  assign N34 = N266;
  assign data_mem_addr_li[53:45] = (N35)? dcache_pkt_i[75:67] : 
                                   (N275)? wbuf_entry_out[86:78] : 
                                   (N271)? { lce_data_mem_pkt[521:516], N272, lce_data_mem_pkt[514:514], N273 } : 1'b0;
  assign N35 = N268;
  assign data_mem_data_li[383:320] = (N36)? wbuf_entry_out[74:11] : 
                                     (N37)? lce_data_mem_write_data[383:320] : 1'b0;
  assign N36 = N277;
  assign N37 = N276;
  assign data_mem_mask_li[47:40] = (N38)? wbuf_entry_out[10:3] : 
                                   (N39)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N38 = N279;
  assign N39 = N278;
  assign data_mem_addr_li[62:54] = (N40)? dcache_pkt_i[75:67] : 
                                   (N287)? wbuf_entry_out[86:78] : 
                                   (N283)? { lce_data_mem_pkt[521:516], N284, N285, lce_data_mem_pkt[513:513] } : 1'b0;
  assign N40 = N280;
  assign data_mem_data_li[447:384] = (N41)? wbuf_entry_out[74:11] : 
                                     (N42)? lce_data_mem_write_data[447:384] : 1'b0;
  assign N41 = N289;
  assign N42 = N288;
  assign data_mem_mask_li[55:48] = (N43)? wbuf_entry_out[10:3] : 
                                   (N44)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N43 = N291;
  assign N44 = N290;
  assign data_mem_addr_li[71:63] = (N45)? dcache_pkt_i[75:67] : 
                                   (N300)? wbuf_entry_out[86:78] : 
                                   (N295)? { lce_data_mem_pkt[521:516], N296, N297, N298 } : 1'b0;
  assign N45 = N292;
  assign data_mem_data_li[511:448] = (N46)? wbuf_entry_out[74:11] : 
                                     (N47)? lce_data_mem_write_data[511:448] : 1'b0;
  assign N46 = N302;
  assign N47 = N301;
  assign data_mem_mask_li[63:56] = (N48)? wbuf_entry_out[10:3] : 
                                   (N49)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N48 = N304;
  assign N49 = N303;
  assign tag_mem_addr_li = (N50)? dcache_pkt_i[75:70] : 
                           (N51)? lce_tag_mem_pkt[22:17] : 1'b0;
  assign N50 = tl_we;
  assign N51 = N472;
  assign tag_mem_data_li = (N52)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N53)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N54)? { lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2] } : 
                           (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N52 = N307;
  assign N53 = N309;
  assign N54 = N311;
  assign N55 = N312;
  assign tag_mem_mask_li = (N52)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                           (N53)? { lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N54)? { lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0] } : 
                           (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_li = (N56)? N314 : 
                         (N57)? N315 : 1'b0;
  assign N56 = v_tv_r;
  assign N57 = N313;
  assign stat_mem_addr_li = (N56)? paddr_tv_r[11:6] : 
                            (N57)? lce_stat_mem_pkt[10:5] : 1'b0;
  assign { N319, N318, N317 } = (N58)? store_hit_way : 
                                (N59)? load_hit_way : 1'b0;
  assign N58 = store_op_tv_r;
  assign N59 = N316;
  assign { N340, N339, N338, N337, N336, N335, N334 } = (N60)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N61)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N62)? { N327, N328, N329, N330, N331, N332, N333 } : 
                                                        (N63)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N60 = N321;
  assign N61 = N323;
  assign N62 = N324;
  assign N63 = N326;
  assign { N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341 } = (N60)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                        (N61)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, dirty_mask_lo } : 
                                                                                                        (N62)? { lru_decode_mask_lo, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                        (N63)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lru_decode_way_li = (N64)? { N319, N318, N317 } : 
                             (N57)? lce_stat_mem_pkt[4:2] : 1'b0;
  assign N64 = stat_mem_data_li[0];
  assign dirty_mask_way_li = (N64)? store_hit_way : 
                             (N57)? lce_stat_mem_pkt[4:2] : 1'b0;
  assign dirty_mask_v_li = (N64)? store_op_tv_r : 
                           (N57)? 1'b1 : 1'b0;
  assign stat_mem_data_li[14:1] = (N64)? { lru_decode_data_lo, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                  (N57)? { N340, N339, N338, N337, N336, N335, N334, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_mask_li = (N64)? { lru_decode_mask_lo, dirty_mask_lo } : 
                            (N57)? { N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341 } : 1'b0;
  assign load_op = ~dcache_pkt_i[79];
  assign signed_op = ~dcache_pkt_i[78];
  assign tl_we = N414 & N415;
  assign N414 = v_i & ready_o;
  assign N415 = ~poison_i;
  assign N65 = ~reset_i;
  assign N66 = reset_i;
  assign N67 = tl_we & dcache_pkt_i[79];
  assign n_0_net_ = N416 & tag_mem_v_li;
  assign N416 = ~reset_i;
  assign n_1_net_ = N417 & data_mem_v_li[0];
  assign N417 = ~reset_i;
  assign n_2_net_ = N418 & data_mem_v_li[1];
  assign N418 = ~reset_i;
  assign n_3_net_ = N419 & data_mem_v_li[2];
  assign N419 = ~reset_i;
  assign n_4_net_ = N420 & data_mem_v_li[3];
  assign N420 = ~reset_i;
  assign n_5_net_ = N421 & data_mem_v_li[4];
  assign N421 = ~reset_i;
  assign n_6_net_ = N422 & data_mem_v_li[5];
  assign N422 = ~reset_i;
  assign n_7_net_ = N423 & data_mem_v_li[6];
  assign N423 = ~reset_i;
  assign n_8_net_ = N424 & data_mem_v_li[7];
  assign N424 = ~reset_i;
  assign tv_we = N425 & N426;
  assign N425 = v_tl_r & N415;
  assign N426 = ~tlb_miss_i;
  assign N71 = ~reset_i;
  assign N72 = reset_i;
  assign N73 = tv_we & load_op_tl_r;
  assign N74 = tv_we & store_op_tl_r;
  assign load_hit_tv[0] = N85 & N380;
  assign store_hit_tv[0] = N86 & N404;
  assign load_hit_tv[1] = N87 & N379;
  assign store_hit_tv[1] = N88 & N401;
  assign load_hit_tv[2] = N89 & N378;
  assign store_hit_tv[2] = N90 & N398;
  assign load_hit_tv[3] = N91 & N377;
  assign store_hit_tv[3] = N92 & N395;
  assign load_hit_tv[4] = N93 & N376;
  assign store_hit_tv[4] = N94 & N392;
  assign load_hit_tv[5] = N95 & N375;
  assign store_hit_tv[5] = N96 & N389;
  assign load_hit_tv[6] = N97 & N374;
  assign store_hit_tv[6] = N98 & N386;
  assign load_hit_tv[7] = N99 & N373;
  assign store_hit_tv[7] = N100 & N383;
  assign load_miss_tv = N428 & load_op_tv_r;
  assign N428 = N427 & v_tv_r;
  assign N427 = ~load_hit;
  assign store_miss_tv = N430 & store_op_tv_r;
  assign N430 = N429 & v_tv_r;
  assign N429 = ~store_hit;
  assign N101 = word_op_tv_r | double_op_tv_r;
  assign N102 = half_op_tv_r | N101;
  assign N103 = ~N102;
  assign N104 = ~double_op_tv_r;
  assign N105 = word_op_tv_r & N104;
  assign N106 = ~word_op_tv_r;
  assign N107 = N104 & N106;
  assign N108 = half_op_tv_r & N107;
  assign N109 = word_op_tv_r | double_op_tv_r;
  assign N110 = half_op_tv_r | N109;
  assign N111 = ~N110;
  assign N112 = ~paddr_tv_r[2];
  assign N113 = ~paddr_tv_r[2];
  assign N114 = ~paddr_tv_r[2];
  assign N115 = ~paddr_tv_r[2];
  assign N116 = paddr_tv_r[2] & paddr_tv_r[1];
  assign N117 = paddr_tv_r[2] & paddr_tv_r[1];
  assign N118 = paddr_tv_r[2] & N431;
  assign N431 = ~paddr_tv_r[1];
  assign N119 = paddr_tv_r[2] & N432;
  assign N432 = ~paddr_tv_r[1];
  assign N120 = N433 & paddr_tv_r[1];
  assign N433 = ~paddr_tv_r[2];
  assign N121 = N434 & paddr_tv_r[1];
  assign N434 = ~paddr_tv_r[2];
  assign N122 = N435 & N436;
  assign N435 = ~paddr_tv_r[2];
  assign N436 = ~paddr_tv_r[1];
  assign N123 = N437 & N438;
  assign N437 = ~paddr_tv_r[2];
  assign N438 = ~paddr_tv_r[1];
  assign N124 = N439 & paddr_tv_r[0];
  assign N439 = paddr_tv_r[2] & paddr_tv_r[1];
  assign N125 = N440 & N441;
  assign N440 = paddr_tv_r[2] & paddr_tv_r[1];
  assign N441 = ~paddr_tv_r[0];
  assign N126 = N443 & paddr_tv_r[0];
  assign N443 = paddr_tv_r[2] & N442;
  assign N442 = ~paddr_tv_r[1];
  assign N127 = N445 & N446;
  assign N445 = paddr_tv_r[2] & N444;
  assign N444 = ~paddr_tv_r[1];
  assign N446 = ~paddr_tv_r[0];
  assign N128 = N448 & paddr_tv_r[0];
  assign N448 = N447 & paddr_tv_r[1];
  assign N447 = ~paddr_tv_r[2];
  assign N129 = N450 & N451;
  assign N450 = N449 & paddr_tv_r[1];
  assign N449 = ~paddr_tv_r[2];
  assign N451 = ~paddr_tv_r[0];
  assign N130 = N454 & paddr_tv_r[0];
  assign N454 = N452 & N453;
  assign N452 = ~paddr_tv_r[2];
  assign N453 = ~paddr_tv_r[1];
  assign N131 = N457 & N458;
  assign N457 = N455 & N456;
  assign N455 = ~paddr_tv_r[2];
  assign N456 = ~paddr_tv_r[1];
  assign N458 = ~paddr_tv_r[0];
  assign N132 = word_op_tv_r & N104;
  assign N133 = N104 & N106;
  assign N134 = half_op_tv_r & N133;
  assign n_10_net_ = N459 & stat_mem_v_li;
  assign N459 = ~reset_i;
  assign N135 = ~invalid_exist;
  assign v_o = N462 & N463;
  assign N462 = v_tv_r & N461;
  assign N461 = ~N460;
  assign N460 = load_miss_tv | store_miss_tv;
  assign N463 = ~reset_i;
  assign n_13_net__2_ = load_hit_way[2] ^ paddr_tv_r[5];
  assign n_13_net__1_ = load_hit_way[1] ^ paddr_tv_r[4];
  assign n_13_net__0_ = load_hit_way[0] ^ paddr_tv_r[3];
  assign genblk4_word_sigext = signed_op_tv_r & genblk4_data_word_selected[31];
  assign genblk4_half_sigext = signed_op_tv_r & genblk4_data_half_selected[15];
  assign genblk4_byte_sigext = signed_op_tv_r & genblk4_data_byte_selected[7];
  assign N136 = ~load_op_tv_r;
  assign N137 = word_op_tv_r | double_op_tv_r;
  assign N138 = half_op_tv_r | N137;
  assign N139 = ~N138;
  assign N204 = word_op_tv_r & N104;
  assign N205 = N104 & N106;
  assign N206 = half_op_tv_r & N205;
  assign n_14_net__2_ = wbuf_entry_out[2] ^ wbuf_entry_out[80];
  assign n_14_net__1_ = wbuf_entry_out[1] ^ wbuf_entry_out[79];
  assign n_14_net__0_ = wbuf_entry_out[0] ^ wbuf_entry_out[78];
  assign N207 = load_op & tl_we;
  assign N208 = wbuf_yumi_li;
  assign N209 = N208 | N207;
  assign N210 = ~N209;
  assign N211 = ~N207;
  assign N212 = N208 & N211;
  assign data_mem_w_li[7] = wbuf_yumi_li | N464;
  assign N464 = lce_data_mem_pkt_yumi_li & lce_data_mem_pkt[0];
  assign data_mem_w_li[6] = wbuf_yumi_li | N465;
  assign N465 = lce_data_mem_pkt_yumi_li & lce_data_mem_pkt[0];
  assign data_mem_w_li[5] = wbuf_yumi_li | N466;
  assign N466 = lce_data_mem_pkt_yumi_li & lce_data_mem_pkt[0];
  assign data_mem_w_li[4] = wbuf_yumi_li | N467;
  assign N467 = lce_data_mem_pkt_yumi_li & lce_data_mem_pkt[0];
  assign data_mem_w_li[3] = wbuf_yumi_li | N468;
  assign N468 = lce_data_mem_pkt_yumi_li & lce_data_mem_pkt[0];
  assign data_mem_w_li[2] = wbuf_yumi_li | N469;
  assign N469 = lce_data_mem_pkt_yumi_li & lce_data_mem_pkt[0];
  assign data_mem_w_li[1] = wbuf_yumi_li | N470;
  assign N470 = lce_data_mem_pkt_yumi_li & lce_data_mem_pkt[0];
  assign data_mem_w_li[0] = wbuf_yumi_li | N471;
  assign N471 = lce_data_mem_pkt_yumi_li & lce_data_mem_pkt[0];
  assign N213 = load_op & tl_we;
  assign N214 = wbuf_yumi_li;
  assign N215 = N214 | N213;
  assign N216 = ~N215;
  assign N217 = ~N213;
  assign N218 = N214 & N217;
  assign N219 = ~wbuf_yumi_li;
  assign N220 = wbuf_yumi_li;
  assign N221 = ~wbuf_yumi_li;
  assign N222 = wbuf_yumi_li;
  assign N223 = load_op & tl_we;
  assign N224 = wbuf_yumi_li;
  assign N225 = N224 | N223;
  assign N226 = ~N225;
  assign N227 = ~lce_data_mem_pkt[513];
  assign N228 = ~N223;
  assign N229 = N224 & N228;
  assign n_18_net__0_ = ~lce_data_mem_pkt[513];
  assign N230 = ~wbuf_yumi_li;
  assign N231 = wbuf_yumi_li;
  assign N232 = ~wbuf_yumi_li;
  assign N233 = wbuf_yumi_li;
  assign N234 = load_op & tl_we;
  assign N235 = wbuf_yumi_li;
  assign N236 = N235 | N234;
  assign N237 = ~N236;
  assign N238 = ~lce_data_mem_pkt[514];
  assign N239 = ~N234;
  assign N240 = N235 & N239;
  assign n_20_net__1_ = ~lce_data_mem_pkt[514];
  assign N241 = ~wbuf_yumi_li;
  assign N242 = wbuf_yumi_li;
  assign N243 = ~wbuf_yumi_li;
  assign N244 = wbuf_yumi_li;
  assign N245 = load_op & tl_we;
  assign N246 = wbuf_yumi_li;
  assign N247 = N246 | N245;
  assign N248 = ~N247;
  assign N249 = ~lce_data_mem_pkt[514];
  assign N250 = ~lce_data_mem_pkt[513];
  assign N251 = ~N245;
  assign N252 = N246 & N251;
  assign n_22_net__1_ = ~lce_data_mem_pkt[514];
  assign n_22_net__0_ = ~lce_data_mem_pkt[513];
  assign N253 = ~wbuf_yumi_li;
  assign N254 = wbuf_yumi_li;
  assign N255 = ~wbuf_yumi_li;
  assign N256 = wbuf_yumi_li;
  assign N257 = load_op & tl_we;
  assign N258 = wbuf_yumi_li;
  assign N259 = N258 | N257;
  assign N260 = ~N259;
  assign N261 = ~lce_data_mem_pkt[515];
  assign N262 = ~N257;
  assign N263 = N258 & N262;
  assign n_24_net__2_ = ~lce_data_mem_pkt[515];
  assign N264 = ~wbuf_yumi_li;
  assign N265 = wbuf_yumi_li;
  assign N266 = ~wbuf_yumi_li;
  assign N267 = wbuf_yumi_li;
  assign N268 = load_op & tl_we;
  assign N269 = wbuf_yumi_li;
  assign N270 = N269 | N268;
  assign N271 = ~N270;
  assign N272 = ~lce_data_mem_pkt[515];
  assign N273 = ~lce_data_mem_pkt[513];
  assign N274 = ~N268;
  assign N275 = N269 & N274;
  assign n_26_net__2_ = ~lce_data_mem_pkt[515];
  assign n_26_net__0_ = ~lce_data_mem_pkt[513];
  assign N276 = ~wbuf_yumi_li;
  assign N277 = wbuf_yumi_li;
  assign N278 = ~wbuf_yumi_li;
  assign N279 = wbuf_yumi_li;
  assign N280 = load_op & tl_we;
  assign N281 = wbuf_yumi_li;
  assign N282 = N281 | N280;
  assign N283 = ~N282;
  assign N284 = ~lce_data_mem_pkt[515];
  assign N285 = ~lce_data_mem_pkt[514];
  assign N286 = ~N280;
  assign N287 = N281 & N286;
  assign n_28_net__2_ = ~lce_data_mem_pkt[515];
  assign n_28_net__1_ = ~lce_data_mem_pkt[514];
  assign N288 = ~wbuf_yumi_li;
  assign N289 = wbuf_yumi_li;
  assign N290 = ~wbuf_yumi_li;
  assign N291 = wbuf_yumi_li;
  assign N292 = load_op & tl_we;
  assign N293 = wbuf_yumi_li;
  assign N294 = N293 | N292;
  assign N295 = ~N294;
  assign N296 = ~lce_data_mem_pkt[515];
  assign N297 = ~lce_data_mem_pkt[514];
  assign N298 = ~lce_data_mem_pkt[513];
  assign N299 = ~N292;
  assign N300 = N293 & N299;
  assign n_30_net__2_ = ~lce_data_mem_pkt[515];
  assign n_30_net__1_ = ~lce_data_mem_pkt[514];
  assign n_30_net__0_ = ~lce_data_mem_pkt[513];
  assign N301 = ~wbuf_yumi_li;
  assign N302 = wbuf_yumi_li;
  assign N303 = ~wbuf_yumi_li;
  assign N304 = wbuf_yumi_li;
  assign tag_mem_v_li = tl_we | lce_tag_mem_pkt_yumi_li;
  assign tag_mem_w_li = N472 & lce_tag_mem_pkt_v_lo;
  assign N472 = ~tl_we;
  assign N305 = ~lce_tag_mem_pkt[1];
  assign N306 = ~lce_tag_mem_pkt[0];
  assign N309 = ~N308;
  assign N311 = ~N310;
  assign stat_mem_v_li = v_tv_r | lce_stat_mem_pkt_yumi_li;
  assign N313 = ~v_tv_r;
  assign N314 = ~N473;
  assign N473 = load_miss_tv | store_miss_tv;
  assign N315 = lce_stat_mem_pkt_yumi_li & N406;
  assign stat_mem_data_li[0] = v_tv_r;
  assign N316 = ~store_op_tv_r;
  assign N320 = ~lce_stat_mem_pkt[1];
  assign N323 = ~N322;
  assign N326 = ~N325;
  assign N327 = ~lru_decode_data_lo[6];
  assign N328 = ~lru_decode_data_lo[5];
  assign N329 = ~lru_decode_data_lo[4];
  assign N330 = ~lru_decode_data_lo[3];
  assign N331 = ~lru_decode_data_lo[2];
  assign N332 = ~lru_decode_data_lo[1];
  assign N333 = ~lru_decode_data_lo[0];
  assign wbuf_v_li = N474 & store_hit;
  assign N474 = v_tv_r & store_op_tv_r;
  assign wbuf_yumi_li = wbuf_v_lo & N476;
  assign N476 = ~N475;
  assign N475 = load_op & tl_we;
  assign bypass_v_li = tv_we & load_op_tl_r;
  assign N356 = N477 & N478;
  assign N477 = lce_data_mem_pkt_v_lo & lce_data_mem_pkt_yumi_li;
  assign N478 = ~lce_data_mem_pkt[0];
  assign n_33_net__0_ = ~lce_data_mem_pkt_way_r[0];
  assign n_34_net__1_ = ~lce_data_mem_pkt_way_r[1];
  assign n_35_net__1_ = ~lce_data_mem_pkt_way_r[1];
  assign n_35_net__0_ = ~lce_data_mem_pkt_way_r[0];
  assign n_36_net__2_ = ~lce_data_mem_pkt_way_r[2];
  assign n_37_net__2_ = ~lce_data_mem_pkt_way_r[2];
  assign n_37_net__0_ = ~lce_data_mem_pkt_way_r[0];
  assign n_38_net__2_ = ~lce_data_mem_pkt_way_r[2];
  assign n_38_net__1_ = ~lce_data_mem_pkt_way_r[1];
  assign n_39_net__2_ = ~lce_data_mem_pkt_way_r[2];
  assign n_39_net__1_ = ~lce_data_mem_pkt_way_r[1];
  assign n_39_net__0_ = ~lce_data_mem_pkt_way_r[0];
  assign lce_data_mem_pkt_yumi_li = N484 & lce_data_mem_pkt_v_lo;
  assign N484 = N482 & N483;
  assign N482 = N480 & N481;
  assign N480 = ~N479;
  assign N479 = load_op & tl_we;
  assign N481 = ~wbuf_v_lo;
  assign N483 = ~lce_snoop_match_lo;
  assign lce_tag_mem_pkt_yumi_li = lce_tag_mem_pkt_v_lo & N472;
  assign lce_stat_mem_pkt_yumi_li = N313 & lce_stat_mem_pkt_v_lo;

  always @(posedge clk_i) begin
    if(N70) begin
      { data_tl_r[63:0] } <= { dcache_pkt_i[63:0] };
    end 
    if(1'b1) begin
      v_tl_r <= N68;
      v_tv_r <= N75;
    end 
    if(N69) begin
      { page_offset_tl_r[11:0] } <= { dcache_pkt_i[75:64] };
      load_op_tl_r <= load_op;
      store_op_tl_r <= dcache_pkt_i[79];
      signed_op_tl_r <= signed_op;
      double_op_tl_r <= N407;
      word_op_tl_r <= N410;
      half_op_tl_r <= N413;
    end 
    if(N84) begin
      { data_tv_r[63:0] } <= { data_tl_r[63:0] };
    end 
    if(N76) begin
      { tag_info_tv_r[95:0] } <= { tag_mem_data_lo[95:0] };
      load_op_tv_r <= load_op_tl_r;
      { paddr_tv_r[21:19] } <= { ptag_i[9:7] };
    end 
    if(N77) begin
      store_op_tv_r <= store_op_tl_r;
      double_op_tv_r <= double_op_tl_r;
      signed_op_tv_r <= signed_op_tl_r;
      word_op_tv_r <= word_op_tl_r;
      half_op_tv_r <= half_op_tl_r;
      { paddr_tv_r[18:0] } <= { ptag_i[6:0], page_offset_tl_r[11:0] };
    end 
    if(N78) begin
      { ld_data_tv_r[511:413], ld_data_tv_r[0:0] } <= { data_mem_data_lo[511:413], data_mem_data_lo[0:0] };
    end 
    if(N79) begin
      { ld_data_tv_r[412:314], ld_data_tv_r[1:1] } <= { data_mem_data_lo[412:314], data_mem_data_lo[1:1] };
    end 
    if(N80) begin
      { ld_data_tv_r[313:215], ld_data_tv_r[2:2] } <= { data_mem_data_lo[313:215], data_mem_data_lo[2:2] };
    end 
    if(N81) begin
      { ld_data_tv_r[214:116], ld_data_tv_r[3:3] } <= { data_mem_data_lo[214:116], data_mem_data_lo[3:3] };
    end 
    if(N82) begin
      { ld_data_tv_r[115:17], ld_data_tv_r[4:4] } <= { data_mem_data_lo[115:17], data_mem_data_lo[4:4] };
    end 
    if(N83) begin
      { ld_data_tv_r[16:5] } <= { data_mem_data_lo[16:5] };
    end 
    if(N356) begin
      { lce_data_mem_pkt_way_r[2:0] } <= { lce_data_mem_pkt[515:513] };
    end 
  end


endmodule



module bp_be_mmu_top_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_num_cce_p1_num_lce_p2_cce_block_size_in_bytes_p64_lce_assoc_p8_lce_sets_p64
(
  clk_i,
  reset_i,
  mmu_cmd_i,
  mmu_cmd_v_i,
  mmu_cmd_ready_o,
  chk_psn_ex_i,
  mmu_resp_o,
  mmu_resp_v_o,
  mmu_resp_ready_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_tr_resp_i,
  lce_tr_resp_v_i,
  lce_tr_resp_ready_o,
  lce_tr_resp_o,
  lce_tr_resp_v_o,
  lce_tr_resp_ready_i,
  dcache_id_i
);

  input [123:0] mmu_cmd_i;
  output [70:0] mmu_resp_o;
  output [29:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [539:0] lce_data_cmd_i;
  input [538:0] lce_tr_resp_i;
  output [538:0] lce_tr_resp_o;
  input [0:0] dcache_id_i;
  input clk_i;
  input reset_i;
  input mmu_cmd_v_i;
  input chk_psn_ex_i;
  input mmu_resp_ready_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_tr_resp_v_i;
  input lce_tr_resp_ready_i;
  output mmu_cmd_ready_o;
  output mmu_resp_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_tr_resp_ready_o;
  output lce_tr_resp_v_o;
  wire [70:0] mmu_resp_o;
  wire [29:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [538:0] lce_tr_resp_o;
  wire mmu_cmd_ready_o,mmu_resp_v_o,lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,
  lce_cmd_ready_o,lce_data_cmd_ready_o,lce_tr_resp_ready_o,lce_tr_resp_v_o,mmu_resp_o_6,
  mmu_resp_o_5,mmu_resp_o_4,mmu_resp_o_3,mmu_resp_o_2,mmu_resp_o_1,dcache_ready,N0;
  reg [9:0] ptag_r;

  bp_be_dcache_data_width_p64_paddr_width_p22_sets_p64_ways_p8_num_cce_p1_num_lce_p2
  dcache
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_id_i(dcache_id_i[0]),
    .dcache_pkt_i({ mmu_cmd_i[123:120], mmu_cmd_i[75:0] }),
    .v_i(mmu_cmd_v_i),
    .ready_o(dcache_ready),
    .data_o(mmu_resp_o[70:7]),
    .v_o(mmu_resp_v_o),
    .tlb_miss_i(1'b0),
    .ptag_i(ptag_r),
    .cache_miss_o(mmu_resp_o[0]),
    .poison_i(chk_psn_ex_i),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_tr_resp_i(lce_tr_resp_i),
    .lce_tr_resp_v_i(lce_tr_resp_v_i),
    .lce_tr_resp_ready_o(lce_tr_resp_ready_o),
    .lce_tr_resp_o(lce_tr_resp_o),
    .lce_tr_resp_v_o(lce_tr_resp_v_o),
    .lce_tr_resp_ready_i(lce_tr_resp_ready_i)
  );

  assign mmu_cmd_ready_o = dcache_ready & N0;
  assign N0 = ~mmu_resp_o[0];

  always @(posedge clk_i) begin
    if(1'b1) begin
      { ptag_r[9:0] } <= { mmu_cmd_i[85:76] };
    end 
  end


endmodule



module bp_be_top
(
  clk_i,
  reset_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_o,
  fe_queue_clr_o,
  fe_queue_dequeue_o,
  fe_queue_rollback_o,
  fe_cmd_o,
  fe_cmd_v_o,
  fe_cmd_ready_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_tr_resp_i,
  lce_tr_resp_v_i,
  lce_tr_resp_ready_o,
  lce_tr_resp_o,
  lce_tr_resp_v_o,
  lce_tr_resp_ready_i,
  proc_cfg_i,
  cmt_trace_stage_reg_o,
  cmt_trace_result_o,
  cmt_trace_exc_o
);

  input [133:0] fe_queue_i;
  output [108:0] fe_cmd_o;
  output [29:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [539:0] lce_data_cmd_i;
  input [538:0] lce_tr_resp_i;
  output [538:0] lce_tr_resp_o;
  input [2:0] proc_cfg_i;
  output [377:0] cmt_trace_stage_reg_o;
  output [127:0] cmt_trace_result_o;
  output [6:0] cmt_trace_exc_o;
  input clk_i;
  input reset_i;
  input fe_queue_v_i;
  input fe_cmd_ready_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_tr_resp_v_i;
  input lce_tr_resp_ready_i;
  output fe_queue_ready_o;
  output fe_queue_clr_o;
  output fe_queue_dequeue_o;
  output fe_queue_rollback_o;
  output fe_cmd_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_tr_resp_ready_o;
  output lce_tr_resp_v_o;
  wire [108:0] fe_cmd_o;
  wire [29:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [538:0] lce_tr_resp_o;
  wire [377:0] cmt_trace_stage_reg_o;
  wire [127:0] cmt_trace_result_o;
  wire [6:0] cmt_trace_exc_o;
  wire fe_queue_ready_o,fe_queue_clr_o,fe_queue_dequeue_o,fe_queue_rollback_o,
  fe_cmd_v_o,lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,
  lce_data_cmd_ready_o,lce_tr_resp_ready_o,lce_tr_resp_v_o,chk_dispatch_v,chk_roll,chk_psn_isd,
  chk_psn_ex,mmu_cmd_rdy,issue_pkt_v,issue_pkt_rdy,mmu_cmd_v,mmu_resp_v,mmu_resp_rdy;
  wire [301:0] calc_status;
  wire [220:0] issue_pkt;
  wire [3:0] decoded_fu_op_n;
  wire [123:0] mmu_cmd;
  wire [70:0] mmu_resp;
  reg [3:0] decoded_fu_op_r;

  bp_be_checker_top_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
  be_checker
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fe_cmd_o(fe_cmd_o),
    .fe_cmd_v_o(fe_cmd_v_o),
    .fe_cmd_ready_i(fe_cmd_ready_i),
    .fe_queue_i(fe_queue_i),
    .fe_queue_v_i(fe_queue_v_i),
    .fe_queue_ready_o(fe_queue_ready_o),
    .chk_roll_fe_o(fe_queue_rollback_o),
    .chk_flush_fe_o(fe_queue_clr_o),
    .chk_dequeue_fe_o(fe_queue_dequeue_o),
    .issue_pkt_o(issue_pkt),
    .issue_pkt_v_o(issue_pkt_v),
    .issue_pkt_ready_i(issue_pkt_rdy),
    .calc_status_i(calc_status),
    .mmu_cmd_ready_i(mmu_cmd_rdy),
    .chk_dispatch_v_o(chk_dispatch_v),
    .chk_roll_o(chk_roll),
    .chk_poison_isd_o(chk_psn_isd),
    .chk_poison_ex_o(chk_psn_ex)
  );


  bp_be_calculator_top_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_core_els_p1_num_lce_p2_lce_sets_p64_cce_block_size_in_bytes_p64
  be_calculator
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .proc_cfg_i(proc_cfg_i),
    .issue_pkt_i(issue_pkt),
    .issue_pkt_v_i(issue_pkt_v),
    .issue_pkt_ready_o(issue_pkt_rdy),
    .chk_dispatch_v_i(chk_dispatch_v),
    .chk_roll_i(chk_roll),
    .chk_poison_ex_i(chk_psn_ex),
    .chk_poison_isd_i(chk_psn_isd),
    .calc_status_o(calc_status),
    .mmu_cmd_o(mmu_cmd),
    .mmu_cmd_v_o(mmu_cmd_v),
    .mmu_cmd_ready_i(mmu_cmd_rdy),
    .mmu_resp_i(mmu_resp),
    .mmu_resp_v_i(mmu_resp_v),
    .mmu_resp_ready_o(mmu_resp_rdy),
    .cmt_trace_stage_reg_o(cmt_trace_stage_reg_o),
    .cmt_trace_result_o(cmt_trace_result_o),
    .cmt_trace_exc_o(cmt_trace_exc_o),
    .decoded_fu_op_o(decoded_fu_op_n)
  );


  bp_be_mmu_top_vaddr_width_p56_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_num_cce_p1_num_lce_p2_cce_block_size_in_bytes_p64_lce_assoc_p8_lce_sets_p64
  be_mmu
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .mmu_cmd_i({ decoded_fu_op_r, mmu_cmd[119:0] }),
    .mmu_cmd_v_i(mmu_cmd_v),
    .mmu_cmd_ready_o(mmu_cmd_rdy),
    .chk_psn_ex_i(chk_psn_ex),
    .mmu_resp_o(mmu_resp),
    .mmu_resp_v_o(mmu_resp_v),
    .mmu_resp_ready_i(mmu_resp_rdy),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_tr_resp_i(lce_tr_resp_i),
    .lce_tr_resp_v_i(lce_tr_resp_v_i),
    .lce_tr_resp_ready_o(lce_tr_resp_ready_o),
    .lce_tr_resp_o(lce_tr_resp_o),
    .lce_tr_resp_v_o(lce_tr_resp_v_o),
    .lce_tr_resp_ready_i(lce_tr_resp_ready_i),
    .dcache_id_i(proc_cfg_i[0])
  );


  always @(posedge clk_i) begin
    if(1'b1) begin
      { decoded_fu_op_r[3:0] } <= { decoded_fu_op_n[3:0] };
    end 
  end


endmodule

