VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO test
  FOREIGN test ;


  SIZE 100.8 BY 100.8 ;
  CLASS BLOCK ;
  PIN in[0]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 19.884999999999998
           98.7
           20.585
           100.8 ;
    END
  END in[0]
  PIN in[1]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 40.025
           98.7
           40.725
           100.8 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 60.165
           98.7
           60.865
           100.8 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 80.305
           98.7
           81.005
           100.8 ;
    END
  END in[3]
  PIN in[12]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 19.884999999999998
           0.0
           20.585
           2.1 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 40.025
           0.0
           40.725
           2.1 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 60.165
           0.0
           60.865
           2.1 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 80.305
           0.0
           81.005
           2.1 ;
    END
  END in[15]
  PIN in[4]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 98.7
           19.74
           100.8
           20.44 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 98.7
           40.04
           100.8
           40.74 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 98.7
           60.06
           100.8
           60.760000000000005 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 98.7
           80.22000000000001
           100.8
           80.92 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.0
           19.74
           2.1
           20.44 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.0
           40.04
           2.1
           40.74 ;
    END
  END in[9]
  PIN in[10]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.0
           60.06
           2.1
           60.760000000000005 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.0
           80.22000000000001
           2.1
           80.92 ;
    END
  END in[11]

  OBS
    LAYER metal1 ;
    RECT 0 0 100.8 100.8 ;
  END
  OBS
    LAYER metal2 ;
    RECT 0 0 100.8 100.8 ;
  END

END test

END LIBRARY