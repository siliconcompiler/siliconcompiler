module or2 (
    input  a,
    input  b,
    output c
);

    assign c = a | b;

endmodule
