(* blackbox *)
module heartbeat (
    input _vdd,
    input _vss,

    input clk,
    input nreset,
    output reg out
);

endmodule
