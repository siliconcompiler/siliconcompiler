# BSD 3-Clause License
# 
# Copyright 2020 Lawrence T. Clark, Vinay Vashishtha, or Arizona State
# University
# 
# Redistribution and use in source and binary forms, with or without
# modification, are permitted provided that the following conditions are met:
# 
# 1. Redistributions of source code must retain the above copyright notice,
# this list of conditions and the following disclaimer.
# 
# 2. Redistributions in binary form must reproduce the above copyright
# notice, this list of conditions and the following disclaimer in the
# documentation and/or other materials provided with the distribution.
# 
# 3. Neither the name of the copyright holder nor the names of its
# contributors may be used to endorse or promote products derived from this
# software without specific prior written permission.
# 
# THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
# AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
# IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
# ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
# LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
# CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
# SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
# INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
# CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
# ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
# POSSIBILITY OF SUCH DAMAGE.

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE asap7sc7p5t
 CLASS CORE ;
 SIZE 0.054 BY 0.270 ;
 SYMMETRY Y ;
END asap7sc7p5t

MACRO A2O1A1Ixp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN A2O1A1Ixp33_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.081 0.252 0.19 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.214 0.215 0.306 0.233 ;
        RECT 0.288 0.037 0.306 0.233 ;
        RECT 0.262 0.037 0.306 0.055 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.23 0.045 ;
      RECT 0.04 0.225 0.176 0.243 ;
  END
END A2O1A1Ixp33_ASAP7_75t_L

MACRO A2O1A1O1Ixp25_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN A2O1A1O1Ixp25_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.127 0.414 0.145 ;
        RECT 0.342 0.07 0.36 0.2 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.261 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.207 0.225 0.387 0.243 ;
      RECT 0.04 0.027 0.225 0.045 ;
      RECT 0.04 0.225 0.171 0.243 ;
  END
END A2O1A1O1Ixp25_ASAP7_75t_L

MACRO AND2x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x2_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.084 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.225 0.306 0.243 ;
        RECT 0.288 0.027 0.306 0.243 ;
        RECT 0.207 0.027 0.306 0.045 ;
        RECT 0.207 0.184 0.225 0.243 ;
        RECT 0.207 0.027 0.225 0.086 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.18 0.243 ;
      RECT 0.162 0.027 0.18 0.243 ;
      RECT 0.162 0.126 0.203 0.144 ;
      RECT 0.07 0.027 0.088 0.086 ;
      RECT 0.07 0.027 0.18 0.045 ;
  END
END AND2x2_ASAP7_75t_L

MACRO AND2x4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x4_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.028 0.252 0.15 ;
        RECT 0.072 0.028 0.252 0.046 ;
        RECT 0.072 0.028 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.107 0.144 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.31 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.231 0.243 ;
      RECT 0.18 0.064 0.198 0.243 ;
      RECT 0.179 0.182 0.306 0.2 ;
      RECT 0.288 0.121 0.306 0.2 ;
      RECT 0.115 0.064 0.198 0.082 ;
  END
END AND2x4_ASAP7_75t_L

MACRO AND2x6_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x6_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.028 0.252 0.15 ;
        RECT 0.072 0.028 0.252 0.046 ;
        RECT 0.072 0.028 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.107 0.144 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.225 0.554 0.243 ;
        RECT 0.31 0.027 0.554 0.045 ;
        RECT 0.45 0.027 0.468 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.231 0.243 ;
      RECT 0.18 0.064 0.198 0.243 ;
      RECT 0.179 0.182 0.306 0.2 ;
      RECT 0.288 0.121 0.306 0.2 ;
      RECT 0.115 0.064 0.198 0.082 ;
  END
END AND2x6_ASAP7_75t_L

MACRO AND3x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x1_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.183 0.306 0.201 ;
        RECT 0.288 0.076 0.306 0.201 ;
        RECT 0.261 0.076 0.306 0.094 ;
        RECT 0.261 0.183 0.279 0.235 ;
        RECT 0.261 0.034 0.279 0.094 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.234 0.243 ;
      RECT 0.216 0.027 0.234 0.243 ;
      RECT 0.216 0.126 0.263 0.144 ;
      RECT 0.04 0.027 0.234 0.045 ;
  END
END AND3x1_ASAP7_75t_L

MACRO AND3x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x2_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.225 0.36 0.243 ;
        RECT 0.342 0.027 0.36 0.243 ;
        RECT 0.261 0.027 0.36 0.045 ;
        RECT 0.261 0.184 0.279 0.243 ;
        RECT 0.261 0.027 0.279 0.086 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.234 0.243 ;
      RECT 0.216 0.027 0.234 0.243 ;
      RECT 0.216 0.126 0.284 0.144 ;
      RECT 0.04 0.027 0.234 0.045 ;
  END
END AND3x2_ASAP7_75t_L

MACRO AND3x4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x4_ASAP7_75t_L 0 0 ;
  SIZE 0.756 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.189 0.649 0.207 ;
        RECT 0.612 0.099 0.649 0.117 ;
        RECT 0.612 0.099 0.63 0.207 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.189 0.541 0.207 ;
        RECT 0.504 0.099 0.541 0.117 ;
        RECT 0.504 0.099 0.522 0.207 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.756 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.23 0.243 ;
        RECT 0.018 0.027 0.23 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.26 0.225 0.746 0.243 ;
      RECT 0.728 0.027 0.746 0.243 ;
      RECT 0.26 0.042 0.278 0.243 ;
      RECT 0.218 0.126 0.278 0.144 ;
      RECT 0.634 0.027 0.746 0.045 ;
      RECT 0.472 0.063 0.701 0.081 ;
      RECT 0.31 0.027 0.554 0.045 ;
  END
END AND3x4_ASAP7_75t_L

MACRO AND4x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x1_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.034 0.198 0.2 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.034 0.252 0.164 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.299 0.225 0.36 0.243 ;
        RECT 0.342 0.027 0.36 0.243 ;
        RECT 0.31 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.225 0.252 0.243 ;
      RECT 0.234 0.189 0.252 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.234 0.189 0.306 0.207 ;
      RECT 0.288 0.12 0.306 0.207 ;
      RECT 0.018 0.027 0.085 0.045 ;
  END
END AND4x1_ASAP7_75t_L

MACRO AND4x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x2_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.034 0.306 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.034 0.252 0.2 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.034 0.198 0.164 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.122 0.243 ;
        RECT 0.018 0.027 0.122 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.153 0.225 0.414 0.243 ;
      RECT 0.396 0.027 0.414 0.243 ;
      RECT 0.153 0.189 0.171 0.243 ;
      RECT 0.099 0.189 0.171 0.207 ;
      RECT 0.099 0.119 0.117 0.207 ;
      RECT 0.364 0.027 0.414 0.045 ;
  END
END AND4x2_ASAP7_75t_L

MACRO AND5x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND5x1_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.034 0.198 0.2 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.034 0.252 0.2 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.034 0.306 0.164 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.349 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.35 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.225 0.306 0.243 ;
      RECT 0.288 0.189 0.306 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.288 0.189 0.36 0.207 ;
      RECT 0.342 0.116 0.36 0.207 ;
      RECT 0.018 0.027 0.07 0.045 ;
  END
END AND5x1_ASAP7_75t_L

MACRO AND5x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND5x2_ASAP7_75t_L 0 0 ;
  SIZE 1.08 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.189 0.757 0.207 ;
        RECT 0.72 0.099 0.757 0.117 ;
        RECT 0.72 0.099 0.738 0.207 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.593 0.189 0.63 0.207 ;
        RECT 0.612 0.099 0.63 0.207 ;
        RECT 0.593 0.099 0.63 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.189 0.487 0.207 ;
        RECT 0.45 0.099 0.487 0.117 ;
        RECT 0.45 0.099 0.468 0.207 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.269 0.189 0.306 0.207 ;
        RECT 0.288 0.099 0.306 0.207 ;
        RECT 0.269 0.099 0.306 0.117 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.08 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.958 0.225 1.062 0.243 ;
        RECT 1.044 0.027 1.062 0.243 ;
        RECT 0.958 0.027 1.062 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.148 0.225 0.9 0.243 ;
      RECT 0.882 0.027 0.9 0.243 ;
      RECT 0.882 0.126 0.942 0.144 ;
      RECT 0.742 0.027 0.9 0.045 ;
      RECT 0.58 0.063 0.824 0.081 ;
      RECT 0.418 0.027 0.662 0.045 ;
      RECT 0.256 0.063 0.5 0.081 ;
      RECT 0.094 0.027 0.338 0.045 ;
  END
END AND5x2_ASAP7_75t_L

MACRO AO211x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211x2_ASAP7_75t_L 0 0 ;
  SIZE 0.864 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.126 0.203 0.144 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.311 0.144 ;
        RECT 0.215 0.189 0.252 0.207 ;
        RECT 0.234 0.063 0.252 0.207 ;
        RECT 0.215 0.063 0.252 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.153 0.541 0.171 ;
        RECT 0.504 0.063 0.522 0.171 ;
        RECT 0.485 0.063 0.522 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.864 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.742 0.225 0.846 0.243 ;
        RECT 0.828 0.027 0.846 0.243 ;
        RECT 0.742 0.027 0.846 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.526 0.225 0.684 0.243 ;
      RECT 0.666 0.027 0.684 0.243 ;
      RECT 0.666 0.125 0.743 0.143 ;
      RECT 0.094 0.027 0.684 0.045 ;
      RECT 0.31 0.189 0.608 0.207 ;
      RECT 0.04 0.225 0.393 0.243 ;
  END
END AO211x2_ASAP7_75t_L

MACRO AO21x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21x1_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.034 0.036 0.207 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.23 0.225 0.295 0.243 ;
        RECT 0.277 0.038 0.295 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.189 0.252 0.207 ;
      RECT 0.234 0.027 0.252 0.207 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.04 0.225 0.176 0.243 ;
  END
END AO21x1_ASAP7_75t_L

MACRO AO21x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21x2_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.034 0.036 0.207 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.23 0.225 0.333 0.243 ;
        RECT 0.315 0.069 0.333 0.243 ;
        RECT 0.276 0.069 0.333 0.087 ;
        RECT 0.276 0.038 0.294 0.087 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.189 0.252 0.207 ;
      RECT 0.234 0.027 0.252 0.207 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.04 0.225 0.176 0.243 ;
  END
END AO21x2_ASAP7_75t_L

MACRO AO221x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221x1_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.225 0.522 0.243 ;
        RECT 0.504 0.027 0.522 0.243 ;
        RECT 0.459 0.027 0.522 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.189 0.126 0.207 ;
      RECT 0.018 0.027 0.036 0.207 ;
      RECT 0.396 0.126 0.474 0.144 ;
      RECT 0.396 0.027 0.414 0.144 ;
      RECT 0.018 0.027 0.414 0.045 ;
      RECT 0.2 0.189 0.339 0.207 ;
      RECT 0.039 0.225 0.176 0.243 ;
  END
END AO221x1_ASAP7_75t_L

MACRO AO221x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221x2_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.225 0.549 0.243 ;
        RECT 0.531 0.027 0.549 0.243 ;
        RECT 0.459 0.027 0.549 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.189 0.126 0.207 ;
      RECT 0.018 0.027 0.036 0.207 ;
      RECT 0.396 0.126 0.474 0.144 ;
      RECT 0.396 0.027 0.414 0.144 ;
      RECT 0.018 0.027 0.414 0.045 ;
      RECT 0.2 0.189 0.339 0.207 ;
      RECT 0.039 0.225 0.176 0.243 ;
  END
END AO221x2_ASAP7_75t_L

MACRO AO222x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222x2_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.2 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.164 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.526 0.225 0.63 0.243 ;
        RECT 0.612 0.027 0.63 0.243 ;
        RECT 0.531 0.027 0.63 0.045 ;
        RECT 0.531 0.027 0.549 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.009 0.189 0.122 0.207 ;
      RECT 0.009 0.027 0.027 0.207 ;
      RECT 0.486 0.126 0.554 0.144 ;
      RECT 0.486 0.027 0.504 0.144 ;
      RECT 0.009 0.027 0.504 0.045 ;
      RECT 0.342 0.225 0.468 0.243 ;
      RECT 0.342 0.189 0.36 0.243 ;
      RECT 0.202 0.189 0.36 0.207 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END AO222x2_ASAP7_75t_L

MACRO AO22x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22x1_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.287 0.081 ;
        RECT 0.234 0.063 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.418 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.189 0.36 0.207 ;
      RECT 0.342 0.027 0.36 0.207 ;
      RECT 0.342 0.126 0.419 0.144 ;
      RECT 0.107 0.027 0.36 0.045 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END AO22x1_ASAP7_75t_L

MACRO AO22x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22x2_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.287 0.081 ;
        RECT 0.234 0.063 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.225 0.522 0.243 ;
        RECT 0.504 0.027 0.522 0.243 ;
        RECT 0.418 0.027 0.522 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.189 0.36 0.207 ;
      RECT 0.342 0.027 0.36 0.207 ;
      RECT 0.342 0.126 0.419 0.144 ;
      RECT 0.107 0.027 0.36 0.045 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END AO22x2_ASAP7_75t_L

MACRO AO31x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31x2_ASAP7_75t_L 0 0 ;
  SIZE 0.864 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.099 0.576 0.149 ;
        RECT 0.504 0.099 0.576 0.117 ;
        RECT 0.485 0.153 0.522 0.171 ;
        RECT 0.504 0.099 0.522 0.171 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.099 0.414 0.149 ;
        RECT 0.288 0.099 0.414 0.117 ;
        RECT 0.288 0.153 0.325 0.171 ;
        RECT 0.288 0.07 0.306 0.171 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.059 0.207 ;
        RECT 0.018 0.027 0.059 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.126 0.203 0.144 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.864 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.225 0.846 0.243 ;
        RECT 0.828 0.027 0.846 0.243 ;
        RECT 0.742 0.027 0.846 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.225 0.684 0.243 ;
      RECT 0.666 0.027 0.684 0.243 ;
      RECT 0.612 0.189 0.63 0.243 ;
      RECT 0.199 0.189 0.63 0.207 ;
      RECT 0.234 0.063 0.252 0.207 ;
      RECT 0.666 0.126 0.797 0.144 ;
      RECT 0.2 0.063 0.252 0.081 ;
      RECT 0.526 0.027 0.684 0.045 ;
      RECT 0.364 0.063 0.608 0.081 ;
      RECT 0.04 0.225 0.554 0.243 ;
      RECT 0.094 0.027 0.447 0.045 ;
  END
END AO31x2_ASAP7_75t_L

MACRO AO322x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO322x2_ASAP7_75t_L 0 0 ;
  SIZE 0.81 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.153 0.325 0.171 ;
        RECT 0.288 0.063 0.325 0.081 ;
        RECT 0.288 0.063 0.306 0.171 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.063 0.541 0.081 ;
        RECT 0.504 0.063 0.522 0.164 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.81 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.634 0.225 0.792 0.243 ;
        RECT 0.774 0.027 0.792 0.243 ;
        RECT 0.634 0.027 0.792 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.189 0.576 0.207 ;
      RECT 0.558 0.126 0.576 0.207 ;
      RECT 0.396 0.027 0.414 0.207 ;
      RECT 0.558 0.126 0.743 0.144 ;
      RECT 0.04 0.027 0.446 0.045 ;
      RECT 0.094 0.225 0.198 0.243 ;
      RECT 0.18 0.189 0.198 0.243 ;
      RECT 0.18 0.189 0.338 0.207 ;
      RECT 0.256 0.225 0.5 0.243 ;
  END
END AO322x2_ASAP7_75t_L

MACRO AO32x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32x1_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.063 0.063 0.081 ;
        RECT 0.045 0.034 0.063 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.31 0.189 0.414 0.207 ;
      RECT 0.396 0.027 0.414 0.207 ;
      RECT 0.062 0.126 0.108 0.144 ;
      RECT 0.09 0.027 0.108 0.144 ;
      RECT 0.09 0.027 0.414 0.045 ;
      RECT 0.148 0.225 0.392 0.243 ;
  END
END AO32x1_ASAP7_75t_L

MACRO AO32x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32x2_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.189 0.33 0.207 ;
        RECT 0.288 0.07 0.306 0.207 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.122 0.243 ;
        RECT 0.018 0.068 0.117 0.086 ;
        RECT 0.099 0.037 0.117 0.086 ;
        RECT 0.018 0.068 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.189 0.468 0.207 ;
      RECT 0.45 0.027 0.468 0.207 ;
      RECT 0.093 0.126 0.162 0.144 ;
      RECT 0.144 0.027 0.162 0.144 ;
      RECT 0.144 0.027 0.468 0.045 ;
      RECT 0.202 0.225 0.446 0.243 ;
  END
END AO32x2_ASAP7_75t_L

MACRO AO331x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO331x1_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.081 0.045 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.471 0.225 0.522 0.243 ;
      RECT 0.504 0.027 0.522 0.243 ;
      RECT 0.072 0.063 0.09 0.152 ;
      RECT 0.072 0.063 0.144 0.081 ;
      RECT 0.126 0.027 0.144 0.081 ;
      RECT 0.126 0.027 0.522 0.045 ;
      RECT 0.308 0.189 0.447 0.207 ;
      RECT 0.146 0.225 0.393 0.243 ;
  END
END AO331x1_ASAP7_75t_L

MACRO AO331x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO331x2_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.07 0.522 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.027 0.135 0.045 ;
        RECT 0.072 0.225 0.122 0.243 ;
        RECT 0.072 0.027 0.09 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.525 0.225 0.576 0.243 ;
      RECT 0.558 0.027 0.576 0.243 ;
      RECT 0.126 0.063 0.144 0.152 ;
      RECT 0.126 0.063 0.198 0.081 ;
      RECT 0.18 0.027 0.198 0.081 ;
      RECT 0.18 0.027 0.576 0.045 ;
      RECT 0.362 0.189 0.501 0.207 ;
      RECT 0.2 0.225 0.447 0.243 ;
  END
END AO331x2_ASAP7_75t_L

MACRO AO332x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO332x1_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.07 0.522 0.164 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.094 0.045 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.471 0.189 0.576 0.207 ;
      RECT 0.558 0.027 0.576 0.207 ;
      RECT 0.072 0.063 0.09 0.151 ;
      RECT 0.072 0.063 0.144 0.081 ;
      RECT 0.126 0.027 0.144 0.081 ;
      RECT 0.126 0.027 0.576 0.045 ;
      RECT 0.146 0.225 0.252 0.243 ;
      RECT 0.234 0.189 0.252 0.243 ;
      RECT 0.234 0.189 0.393 0.207 ;
      RECT 0.308 0.225 0.556 0.243 ;
  END
END AO332x1_ASAP7_75t_L

MACRO AO332x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO332x2_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.07 0.576 0.164 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.07 0.522 0.164 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.148 0.045 ;
        RECT 0.018 0.225 0.122 0.243 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.525 0.189 0.63 0.207 ;
      RECT 0.612 0.027 0.63 0.207 ;
      RECT 0.126 0.063 0.144 0.151 ;
      RECT 0.126 0.063 0.198 0.081 ;
      RECT 0.18 0.027 0.198 0.081 ;
      RECT 0.18 0.027 0.63 0.045 ;
      RECT 0.2 0.225 0.306 0.243 ;
      RECT 0.288 0.189 0.306 0.243 ;
      RECT 0.288 0.189 0.447 0.207 ;
      RECT 0.362 0.225 0.61 0.243 ;
  END
END AO332x2_ASAP7_75t_L

MACRO AO333x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO333x1_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.07 0.576 0.164 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.07 0.522 0.164 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.081 0.045 ;
        RECT 0.018 0.225 0.069 0.243 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.471 0.225 0.63 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.072 0.063 0.09 0.152 ;
      RECT 0.072 0.063 0.144 0.081 ;
      RECT 0.126 0.027 0.144 0.081 ;
      RECT 0.126 0.027 0.63 0.045 ;
      RECT 0.31 0.189 0.576 0.207 ;
      RECT 0.148 0.225 0.395 0.243 ;
  END
END AO333x1_ASAP7_75t_L

MACRO AO333x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO333x2_ASAP7_75t_L 0 0 ;
  SIZE 0.702 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.07 0.63 0.164 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.07 0.576 0.164 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.07 0.522 0.164 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.702 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.122 0.243 ;
        RECT 0.018 0.081 0.117 0.099 ;
        RECT 0.099 0.045 0.117 0.099 ;
        RECT 0.018 0.081 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.525 0.225 0.684 0.243 ;
      RECT 0.666 0.027 0.684 0.243 ;
      RECT 0.067 0.126 0.162 0.144 ;
      RECT 0.144 0.027 0.162 0.144 ;
      RECT 0.144 0.027 0.684 0.045 ;
      RECT 0.364 0.189 0.63 0.207 ;
      RECT 0.202 0.225 0.449 0.243 ;
  END
END AO333x2_ASAP7_75t_L

MACRO AO33x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO33x2_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.122 0.243 ;
        RECT 0.018 0.068 0.117 0.086 ;
        RECT 0.099 0.037 0.117 0.086 ;
        RECT 0.018 0.068 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.361 0.189 0.522 0.207 ;
      RECT 0.504 0.027 0.522 0.207 ;
      RECT 0.067 0.126 0.162 0.144 ;
      RECT 0.144 0.027 0.162 0.144 ;
      RECT 0.144 0.027 0.522 0.045 ;
      RECT 0.199 0.225 0.449 0.243 ;
  END
END AO33x2_ASAP7_75t_L

MACRO AOI211x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211x1_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.126 0.229 0.144 ;
        RECT 0.18 0.189 0.223 0.207 ;
        RECT 0.18 0.063 0.22 0.081 ;
        RECT 0.18 0.063 0.198 0.207 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.123 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.153 0.442 0.171 ;
        RECT 0.396 0.063 0.442 0.081 ;
        RECT 0.396 0.063 0.414 0.171 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.126 0.554 0.144 ;
        RECT 0.504 0.063 0.55 0.081 ;
        RECT 0.504 0.063 0.522 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.519 0.189 0.63 0.207 ;
        RECT 0.612 0.027 0.63 0.207 ;
        RECT 0.091 0.027 0.63 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.091 0.225 0.306 0.243 ;
      RECT 0.288 0.189 0.306 0.243 ;
      RECT 0.288 0.189 0.449 0.207 ;
      RECT 0.361 0.225 0.608 0.243 ;
  END
END AOI211x1_ASAP7_75t_L

MACRO AOI211xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.09 0.144 ;
        RECT 0.018 0.07 0.036 0.2 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.189 0.306 0.207 ;
        RECT 0.288 0.027 0.306 0.207 ;
        RECT 0.04 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.176 0.243 ;
  END
END AOI211xp5_ASAP7_75t_L

MACRO AOI21x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21x1_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.063 0.306 0.164 ;
        RECT 0.126 0.063 0.306 0.081 ;
        RECT 0.126 0.063 0.144 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.19 0.125 0.256 0.143 ;
        RECT 0.19 0.099 0.227 0.171 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.189 0.36 0.207 ;
        RECT 0.342 0.116 0.36 0.207 ;
        RECT 0.072 0.07 0.09 0.207 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.369 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.018 0.027 0.414 0.045 ;
        RECT 0.018 0.225 0.063 0.243 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.225 0.333 0.243 ;
  END
END AOI21x1_ASAP7_75t_L

MACRO AOI21xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.27 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.125 0.095 0.143 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.27 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.225 0.252 0.243 ;
        RECT 0.234 0.027 0.252 0.243 ;
        RECT 0.107 0.027 0.252 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.171 0.243 ;
  END
END AOI21xp33_ASAP7_75t_L

MACRO AOI21xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.27 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.125 0.095 0.143 ;
        RECT 0.018 0.034 0.036 0.2 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.27 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.225 0.252 0.243 ;
        RECT 0.234 0.027 0.252 0.243 ;
        RECT 0.142 0.027 0.252 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.171 0.243 ;
  END
END AOI21xp5_ASAP7_75t_L

MACRO AOI221x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221x1_ASAP7_75t_L 0 0 ;
  SIZE 0.756 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.153 0.217 0.171 ;
        RECT 0.18 0.027 0.198 0.171 ;
        RECT 0.161 0.027 0.198 0.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.126 0.149 0.144 ;
        RECT 0.053 0.153 0.09 0.171 ;
        RECT 0.072 0.027 0.09 0.171 ;
        RECT 0.053 0.027 0.09 0.045 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.081 0.325 0.099 ;
        RECT 0.269 0.153 0.306 0.171 ;
        RECT 0.288 0.081 0.306 0.171 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.153 0.487 0.171 ;
        RECT 0.45 0.081 0.468 0.171 ;
        RECT 0.391 0.126 0.468 0.144 ;
        RECT 0.431 0.081 0.468 0.099 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.126 0.636 0.144 ;
        RECT 0.539 0.189 0.576 0.207 ;
        RECT 0.558 0.081 0.576 0.207 ;
        RECT 0.539 0.081 0.576 0.099 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.756 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.634 0.189 0.738 0.207 ;
        RECT 0.72 0.045 0.738 0.207 ;
        RECT 0.256 0.045 0.738 0.063 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.31 0.225 0.716 0.243 ;
      RECT 0.04 0.189 0.5 0.207 ;
  END
END AOI221x1_ASAP7_75t_L

MACRO AOI221xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.034 0.306 0.164 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.23 0.045 ;
        RECT 0.018 0.189 0.123 0.207 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.201 0.189 0.339 0.207 ;
      RECT 0.04 0.225 0.176 0.243 ;
  END
END AOI221xp5_ASAP7_75t_L

MACRO AOI222xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.034 0.468 0.2 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.399 0.045 ;
        RECT 0.018 0.189 0.122 0.207 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.342 0.225 0.468 0.243 ;
      RECT 0.342 0.189 0.36 0.243 ;
      RECT 0.202 0.189 0.36 0.207 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END AOI222xp33_ASAP7_75t_L

MACRO AOI22x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22x1_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.153 0.379 0.171 ;
        RECT 0.342 0.099 0.379 0.117 ;
        RECT 0.342 0.099 0.36 0.171 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.431 0.153 0.468 0.171 ;
        RECT 0.45 0.063 0.468 0.171 ;
        RECT 0.288 0.063 0.468 0.081 ;
        RECT 0.288 0.063 0.306 0.152 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.161 0.189 0.198 0.207 ;
        RECT 0.18 0.099 0.198 0.207 ;
        RECT 0.161 0.099 0.198 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.252 0.154 ;
        RECT 0.072 0.063 0.252 0.081 ;
        RECT 0.072 0.189 0.109 0.207 ;
        RECT 0.072 0.063 0.09 0.207 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.309 0.189 0.522 0.207 ;
        RECT 0.504 0.027 0.522 0.207 ;
        RECT 0.038 0.027 0.522 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.5 0.243 ;
  END
END AOI22x1_ASAP7_75t_L

MACRO AOI22xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.034 0.09 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.189 0.306 0.207 ;
        RECT 0.288 0.027 0.306 0.207 ;
        RECT 0.148 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END AOI22xp33_ASAP7_75t_L

MACRO AOI22xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.07 0.144 0.207 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.189 0.306 0.207 ;
        RECT 0.288 0.027 0.306 0.207 ;
        RECT 0.148 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END AOI22xp5_ASAP7_75t_L

MACRO AOI311xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI311xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.225 0.36 0.243 ;
        RECT 0.342 0.027 0.36 0.243 ;
        RECT 0.198 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.234 0.243 ;
  END
END AOI311xp33_ASAP7_75t_L

MACRO AOI31xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.034 0.09 0.2 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.189 0.306 0.207 ;
        RECT 0.288 0.027 0.306 0.207 ;
        RECT 0.201 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.093 0.225 0.23 0.243 ;
  END
END AOI31xp33_ASAP7_75t_L

MACRO AOI31xp67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31xp67_ASAP7_75t_L 0 0 ;
  SIZE 0.702 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.666 0.07 0.684 0.2 ;
        RECT 0.553 0.126 0.684 0.144 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.126 0.419 0.144 ;
        RECT 0.288 0.063 0.325 0.081 ;
        RECT 0.288 0.063 0.306 0.164 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.059 0.207 ;
        RECT 0.018 0.027 0.059 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.126 0.203 0.144 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.702 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.585 0.225 0.663 0.243 ;
        RECT 0.585 0.189 0.603 0.243 ;
        RECT 0.202 0.189 0.603 0.207 ;
        RECT 0.234 0.063 0.252 0.207 ;
        RECT 0.202 0.063 0.252 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.526 0.027 0.663 0.045 ;
      RECT 0.364 0.081 0.608 0.099 ;
      RECT 0.04 0.225 0.554 0.243 ;
      RECT 0.094 0.027 0.447 0.045 ;
  END
END AOI31xp67_ASAP7_75t_L

MACRO AOI321xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI321xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.164 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.189 0.414 0.207 ;
        RECT 0.396 0.027 0.414 0.207 ;
        RECT 0.198 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.256 0.225 0.396 0.243 ;
      RECT 0.094 0.189 0.23 0.207 ;
  END
END AOI321xp33_ASAP7_75t_L

MACRO AOI322xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI322xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.165 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.034 0.09 0.164 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.165 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.189 0.468 0.207 ;
        RECT 0.45 0.027 0.468 0.207 ;
        RECT 0.147 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.225 0.45 0.243 ;
      RECT 0.039 0.189 0.284 0.207 ;
  END
END AOI322xp5_ASAP7_75t_L

MACRO AOI32xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.058 0.243 ;
        RECT 0.018 0.063 0.058 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.104 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.104 0.063 0.144 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.189 0.222 0.207 ;
        RECT 0.18 0.07 0.198 0.207 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.189 0.36 0.207 ;
        RECT 0.342 0.027 0.36 0.207 ;
        RECT 0.04 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.338 0.243 ;
  END
END AOI32xp33_ASAP7_75t_L

MACRO AOI331xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI331xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.034 0.09 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.417 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.201 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.254 0.189 0.393 0.207 ;
      RECT 0.092 0.225 0.339 0.243 ;
  END
END AOI331xp33_ASAP7_75t_L

MACRO AOI332xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI332xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.164 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.034 0.09 0.164 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.417 0.189 0.522 0.207 ;
        RECT 0.504 0.027 0.522 0.207 ;
        RECT 0.201 0.027 0.522 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.254 0.225 0.502 0.243 ;
      RECT 0.092 0.189 0.339 0.207 ;
  END
END AOI332xp33_ASAP7_75t_L

MACRO AOI333xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI333xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.07 0.522 0.164 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.164 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.164 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.164 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.034 0.09 0.164 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.413 0.189 0.576 0.207 ;
        RECT 0.558 0.027 0.576 0.207 ;
        RECT 0.201 0.027 0.576 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.254 0.225 0.515 0.243 ;
      RECT 0.094 0.189 0.34 0.207 ;
  END
END AOI333xp33_ASAP7_75t_L

MACRO AOI33xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.034 0.09 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.164 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.189 0.414 0.207 ;
        RECT 0.396 0.027 0.414 0.207 ;
        RECT 0.201 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.225 0.338 0.243 ;
  END
END AOI33xp33_ASAP7_75t_L

MACRO ASYNC_DFFHx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ASYNC_DFFHx1_ASAP7_75t_L 0 0 ;
  SIZE 1.404 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.182 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.088 ;
        RECT 0.099 0.034 0.117 0.088 ;
        RECT 0.072 0.182 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.336 0.225 1.386 0.243 ;
        RECT 1.368 0.027 1.386 0.243 ;
        RECT 1.336 0.027 1.386 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.404 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
    END
  END VSS
  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.632 0.108 1.067 0.126 ;
      LAYER M1 ;
        RECT 1.044 0.103 1.062 0.168 ;
        RECT 0.612 0.18 0.668 0.198 ;
        RECT 0.612 0.108 0.662 0.126 ;
        RECT 0.612 0.108 0.63 0.198 ;
      LAYER V1 ;
        RECT 0.637 0.108 0.655 0.126 ;
        RECT 1.044 0.108 1.062 0.126 ;
    END
  END RESET
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.783 0.072 1.067 0.09 ;
      LAYER M1 ;
        RECT 0.774 0.072 0.811 0.09 ;
        RECT 0.774 0.072 0.792 0.173 ;
      LAYER V1 ;
        RECT 0.788 0.072 0.806 0.09 ;
    END
  END SET
  OBS
    LAYER M1 ;
      RECT 0.963 0.216 1.008 0.234 ;
      RECT 0.963 0.036 0.981 0.234 ;
      RECT 0.918 0.03 0.936 0.217 ;
      RECT 0.858 0.03 0.936 0.048 ;
      RECT 0.558 0.216 0.77 0.234 ;
      RECT 0.693 0.058 0.711 0.234 ;
      RECT 0.558 0.164 0.576 0.234 ;
      RECT 0.418 0.225 0.504 0.243 ;
      RECT 0.486 0.072 0.504 0.243 ;
      RECT 0.486 0.072 0.547 0.09 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.144 0.047 0.162 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.314 0.09 1.332 0.167 ;
      RECT 1.17 0.036 1.202 0.054 ;
      RECT 1.098 0.103 1.116 0.168 ;
      RECT 0.882 0.097 0.9 0.203 ;
      RECT 0.829 0.099 0.847 0.167 ;
      RECT 0.778 0.036 0.819 0.054 ;
      RECT 0.729 0.067 0.747 0.133 ;
      RECT 0.415 0.027 0.608 0.045 ;
      RECT 0.45 0.119 0.468 0.167 ;
      RECT 0.396 0.12 0.414 0.203 ;
      RECT 0.369 0.054 0.387 0.101 ;
      RECT 0.342 0.12 0.36 0.167 ;
      RECT 0.142 0.106 0.16 0.167 ;
    LAYER M2 ;
      RECT 0.913 0.144 1.337 0.162 ;
      RECT 0.783 0.036 1.198 0.054 ;
      RECT 0.741 0.216 1.008 0.234 ;
      RECT 0.175 0.18 0.926 0.198 ;
      RECT 0.019 0.144 0.852 0.162 ;
      RECT 0.364 0.072 0.752 0.09 ;
    LAYER V1 ;
      RECT 1.314 0.144 1.332 0.162 ;
      RECT 1.175 0.036 1.193 0.054 ;
      RECT 1.098 0.144 1.116 0.162 ;
      RECT 0.985 0.216 1.003 0.234 ;
      RECT 0.918 0.144 0.936 0.162 ;
      RECT 0.882 0.18 0.9 0.198 ;
      RECT 0.829 0.144 0.847 0.162 ;
      RECT 0.788 0.036 0.806 0.054 ;
      RECT 0.746 0.216 0.764 0.234 ;
      RECT 0.729 0.072 0.747 0.09 ;
      RECT 0.512 0.072 0.53 0.09 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.396 0.18 0.414 0.198 ;
      RECT 0.369 0.072 0.387 0.09 ;
      RECT 0.342 0.144 0.36 0.162 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END ASYNC_DFFHx1_ASAP7_75t_L

MACRO BUFx10_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx10_ASAP7_75t_L 0 0 ;
  SIZE 0.756 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.756 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.199 0.225 0.738 0.243 ;
        RECT 0.72 0.027 0.738 0.243 ;
        RECT 0.199 0.027 0.738 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.091 0.225 0.144 0.243 ;
      RECT 0.126 0.027 0.144 0.243 ;
      RECT 0.126 0.126 0.689 0.144 ;
      RECT 0.091 0.027 0.144 0.045 ;
  END
END BUFx10_ASAP7_75t_L

MACRO BUFx12_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx12_ASAP7_75t_L 0 0 ;
  SIZE 0.864 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.864 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.199 0.225 0.846 0.243 ;
        RECT 0.828 0.027 0.846 0.243 ;
        RECT 0.199 0.027 0.846 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.144 0.243 ;
      RECT 0.126 0.027 0.144 0.243 ;
      RECT 0.126 0.126 0.8 0.144 ;
      RECT 0.094 0.027 0.144 0.045 ;
  END
END BUFx12_ASAP7_75t_L

MACRO BUFx12f_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx12f_ASAP7_75t_L 0 0 ;
  SIZE 0.972 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.074 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.972 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.972 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.225 0.954 0.243 ;
        RECT 0.936 0.027 0.954 0.243 ;
        RECT 0.31 0.027 0.954 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.279 0.243 ;
      RECT 0.261 0.027 0.279 0.243 ;
      RECT 0.261 0.126 0.311 0.144 ;
      RECT 0.094 0.027 0.279 0.045 ;
  END
END BUFx12f_ASAP7_75t_L

MACRO BUFx16f_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx16f_ASAP7_75t_L 0 0 ;
  SIZE 1.188 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.06 0.243 ;
        RECT 0.018 0.027 0.06 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.225 1.17 0.243 ;
        RECT 1.152 0.027 1.17 0.243 ;
        RECT 0.31 0.027 1.17 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.234 0.126 1.124 0.144 ;
      RECT 0.094 0.027 0.252 0.045 ;
  END
END BUFx16f_ASAP7_75t_L

MACRO BUFx24_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx24_ASAP7_75t_L 0 0 ;
  SIZE 1.62 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.62 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.62 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.225 1.602 0.243 ;
        RECT 1.584 0.027 1.602 0.243 ;
        RECT 0.31 0.027 1.602 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.234 0.126 1.553 0.144 ;
      RECT 0.094 0.027 0.252 0.045 ;
  END
END BUFx24_ASAP7_75t_L

MACRO BUFx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx2_ASAP7_75t_L 0 0 ;
  SIZE 0.27 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.073 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.207 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.27 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.225 0.252 0.243 ;
        RECT 0.234 0.027 0.252 0.243 ;
        RECT 0.145 0.027 0.252 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.12 0.243 ;
      RECT 0.102 0.027 0.12 0.243 ;
      RECT 0.102 0.126 0.203 0.144 ;
      RECT 0.04 0.027 0.12 0.045 ;
  END
END BUFx2_ASAP7_75t_L

MACRO BUFx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx3_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.073 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.207 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.225 0.306 0.243 ;
        RECT 0.288 0.027 0.306 0.243 ;
        RECT 0.145 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.12 0.243 ;
      RECT 0.102 0.027 0.12 0.243 ;
      RECT 0.102 0.126 0.26 0.144 ;
      RECT 0.04 0.027 0.12 0.045 ;
  END
END BUFx3_ASAP7_75t_L

MACRO BUFx4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.073 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.207 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.225 0.357 0.243 ;
        RECT 0.339 0.027 0.357 0.243 ;
        RECT 0.145 0.027 0.357 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.12 0.243 ;
      RECT 0.102 0.027 0.12 0.243 ;
      RECT 0.102 0.126 0.314 0.144 ;
      RECT 0.04 0.027 0.12 0.045 ;
  END
END BUFx4_ASAP7_75t_L

MACRO BUFx4f_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4f_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.098 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.199 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.199 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.091 0.225 0.144 0.243 ;
      RECT 0.126 0.027 0.144 0.243 ;
      RECT 0.126 0.126 0.367 0.144 ;
      RECT 0.091 0.027 0.144 0.045 ;
  END
END BUFx4f_ASAP7_75t_L

MACRO BUFx5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx5_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.073 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.207 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.145 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.12 0.243 ;
      RECT 0.102 0.027 0.12 0.243 ;
      RECT 0.102 0.126 0.368 0.144 ;
      RECT 0.04 0.027 0.12 0.045 ;
  END
END BUFx5_ASAP7_75t_L

MACRO BUFx6f_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx6f_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.084 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.225 0.522 0.243 ;
        RECT 0.504 0.027 0.522 0.243 ;
        RECT 0.202 0.027 0.522 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.144 0.243 ;
      RECT 0.126 0.027 0.144 0.243 ;
      RECT 0.126 0.126 0.473 0.144 ;
      RECT 0.094 0.027 0.144 0.045 ;
  END
END BUFx6f_ASAP7_75t_L

MACRO BUFx8_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx8_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.098 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.225 0.63 0.243 ;
        RECT 0.612 0.027 0.63 0.243 ;
        RECT 0.202 0.027 0.63 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.091 0.225 0.144 0.243 ;
      RECT 0.126 0.027 0.144 0.243 ;
      RECT 0.126 0.126 0.581 0.144 ;
      RECT 0.091 0.027 0.144 0.045 ;
  END
END BUFx8_ASAP7_75t_L

MACRO CKINVDCx10_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx10_ASAP7_75t_L 0 0 ;
  SIZE 1.296 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.088 0.126 1.17 0.144 ;
        RECT 1.12 0.027 1.138 0.144 ;
        RECT 0.05 0.027 1.138 0.045 ;
        RECT 0.764 0.126 0.814 0.144 ;
        RECT 0.796 0.027 0.814 0.144 ;
        RECT 0.374 0.126 0.424 0.144 ;
        RECT 0.374 0.027 0.392 0.144 ;
        RECT 0.05 0.126 0.1 0.144 ;
        RECT 0.05 0.027 0.068 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.296 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.296 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 1.224 0.243 ;
        RECT 1.206 0.063 1.224 0.243 ;
        RECT 1.174 0.063 1.224 0.081 ;
        RECT 1.044 0.063 1.094 0.081 ;
        RECT 1.044 0.063 1.062 0.243 ;
        RECT 0.72 0.063 0.77 0.081 ;
        RECT 0.72 0.063 0.738 0.243 ;
        RECT 0.45 0.063 0.468 0.243 ;
        RECT 0.418 0.063 0.468 0.081 ;
        RECT 0.126 0.063 0.144 0.243 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.936 0.126 0.992 0.144 ;
      RECT 0.936 0.09 0.954 0.144 ;
      RECT 0.85 0.09 1.002 0.108 ;
      RECT 0.831 0.162 0.986 0.18 ;
      RECT 0.882 0.126 0.9 0.18 ;
      RECT 0.842 0.126 0.9 0.144 ;
      RECT 0.526 0.162 0.681 0.18 ;
      RECT 0.612 0.126 0.63 0.18 ;
      RECT 0.612 0.126 0.67 0.144 ;
      RECT 0.52 0.126 0.576 0.144 ;
      RECT 0.558 0.09 0.576 0.144 ;
      RECT 0.51 0.09 0.662 0.108 ;
      RECT 0.202 0.162 0.357 0.18 ;
      RECT 0.288 0.126 0.306 0.18 ;
      RECT 0.288 0.126 0.346 0.144 ;
      RECT 0.196 0.126 0.252 0.144 ;
      RECT 0.234 0.09 0.252 0.144 ;
      RECT 0.186 0.09 0.338 0.108 ;
  END
END CKINVDCx10_ASAP7_75t_L

MACRO CKINVDCx11_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx11_ASAP7_75t_L 0 0 ;
  SIZE 1.404 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.304 0.126 1.354 0.144 ;
        RECT 1.336 0.027 1.354 0.144 ;
        RECT 0.05 0.027 1.354 0.045 ;
        RECT 0.872 0.126 0.964 0.144 ;
        RECT 0.909 0.027 0.927 0.144 ;
        RECT 0.439 0.126 0.531 0.144 ;
        RECT 0.476 0.027 0.494 0.144 ;
        RECT 0.05 0.126 0.1 0.144 ;
        RECT 0.05 0.027 0.068 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.404 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 1.31 0.243 ;
        RECT 1.26 0.063 1.31 0.081 ;
        RECT 1.26 0.063 1.278 0.243 ;
        RECT 0.99 0.063 1.008 0.243 ;
        RECT 0.958 0.063 1.008 0.081 ;
        RECT 0.828 0.063 0.878 0.081 ;
        RECT 0.828 0.063 0.846 0.243 ;
        RECT 0.558 0.063 0.576 0.243 ;
        RECT 0.526 0.063 0.576 0.081 ;
        RECT 0.396 0.063 0.446 0.081 ;
        RECT 0.396 0.063 0.414 0.243 ;
        RECT 0.126 0.063 0.144 0.243 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.152 0.126 1.208 0.144 ;
      RECT 1.152 0.09 1.17 0.144 ;
      RECT 1.066 0.09 1.218 0.108 ;
      RECT 1.047 0.162 1.202 0.18 ;
      RECT 1.098 0.126 1.116 0.18 ;
      RECT 1.058 0.126 1.116 0.144 ;
      RECT 0.634 0.162 0.789 0.18 ;
      RECT 0.72 0.126 0.738 0.18 ;
      RECT 0.72 0.126 0.778 0.144 ;
      RECT 0.628 0.126 0.684 0.144 ;
      RECT 0.666 0.09 0.684 0.144 ;
      RECT 0.618 0.09 0.77 0.108 ;
      RECT 0.202 0.162 0.357 0.18 ;
      RECT 0.288 0.126 0.306 0.18 ;
      RECT 0.288 0.126 0.346 0.144 ;
      RECT 0.196 0.126 0.252 0.144 ;
      RECT 0.234 0.09 0.252 0.144 ;
      RECT 0.186 0.09 0.338 0.108 ;
  END
END CKINVDCx11_ASAP7_75t_L

MACRO CKINVDCx12_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx12_ASAP7_75t_L 0 0 ;
  SIZE 1.404 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.304 0.126 1.354 0.144 ;
        RECT 1.336 0.027 1.354 0.144 ;
        RECT 0.05 0.027 1.354 0.045 ;
        RECT 0.872 0.126 0.964 0.144 ;
        RECT 0.909 0.027 0.927 0.144 ;
        RECT 0.439 0.126 0.531 0.144 ;
        RECT 0.476 0.027 0.494 0.144 ;
        RECT 0.05 0.126 0.1 0.144 ;
        RECT 0.05 0.027 0.068 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.404 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 1.31 0.243 ;
        RECT 1.26 0.063 1.31 0.081 ;
        RECT 1.26 0.063 1.278 0.243 ;
        RECT 0.99 0.063 1.008 0.243 ;
        RECT 0.958 0.063 1.008 0.081 ;
        RECT 0.828 0.063 0.878 0.081 ;
        RECT 0.828 0.063 0.846 0.243 ;
        RECT 0.558 0.063 0.576 0.243 ;
        RECT 0.526 0.063 0.576 0.081 ;
        RECT 0.396 0.063 0.446 0.081 ;
        RECT 0.396 0.063 0.414 0.243 ;
        RECT 0.126 0.063 0.144 0.243 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.152 0.126 1.208 0.144 ;
      RECT 1.152 0.09 1.17 0.144 ;
      RECT 1.066 0.09 1.218 0.108 ;
      RECT 1.047 0.162 1.202 0.18 ;
      RECT 1.098 0.126 1.116 0.18 ;
      RECT 1.058 0.126 1.116 0.144 ;
      RECT 0.634 0.162 0.789 0.18 ;
      RECT 0.72 0.126 0.738 0.18 ;
      RECT 0.72 0.126 0.778 0.144 ;
      RECT 0.628 0.126 0.684 0.144 ;
      RECT 0.666 0.09 0.684 0.144 ;
      RECT 0.618 0.09 0.77 0.108 ;
      RECT 0.202 0.162 0.357 0.18 ;
      RECT 0.288 0.126 0.306 0.18 ;
      RECT 0.288 0.126 0.346 0.144 ;
      RECT 0.196 0.126 0.252 0.144 ;
      RECT 0.234 0.09 0.252 0.144 ;
      RECT 0.186 0.09 0.338 0.108 ;
  END
END CKINVDCx12_ASAP7_75t_L

MACRO CKINVDCx14_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx14_ASAP7_75t_L 0 0 ;
  SIZE 1.512 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.304 0.126 1.397 0.144 ;
        RECT 1.336 0.027 1.354 0.144 ;
        RECT 0.05 0.027 1.354 0.045 ;
        RECT 0.872 0.126 0.964 0.144 ;
        RECT 0.909 0.027 0.927 0.144 ;
        RECT 0.439 0.126 0.531 0.144 ;
        RECT 0.476 0.027 0.494 0.144 ;
        RECT 0.05 0.126 0.1 0.144 ;
        RECT 0.05 0.027 0.068 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.512 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.512 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 1.44 0.243 ;
        RECT 1.422 0.063 1.44 0.243 ;
        RECT 1.39 0.063 1.44 0.081 ;
        RECT 1.26 0.063 1.31 0.081 ;
        RECT 1.26 0.063 1.278 0.243 ;
        RECT 0.99 0.063 1.008 0.243 ;
        RECT 0.958 0.063 1.008 0.081 ;
        RECT 0.828 0.063 0.878 0.081 ;
        RECT 0.828 0.063 0.846 0.243 ;
        RECT 0.558 0.063 0.576 0.243 ;
        RECT 0.526 0.063 0.576 0.081 ;
        RECT 0.396 0.063 0.446 0.081 ;
        RECT 0.396 0.063 0.414 0.243 ;
        RECT 0.126 0.063 0.144 0.243 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.152 0.126 1.208 0.144 ;
      RECT 1.152 0.09 1.17 0.144 ;
      RECT 1.066 0.09 1.218 0.108 ;
      RECT 1.047 0.162 1.202 0.18 ;
      RECT 1.098 0.126 1.116 0.18 ;
      RECT 1.058 0.126 1.116 0.144 ;
      RECT 0.634 0.162 0.789 0.18 ;
      RECT 0.72 0.126 0.738 0.18 ;
      RECT 0.72 0.126 0.778 0.144 ;
      RECT 0.628 0.126 0.684 0.144 ;
      RECT 0.666 0.09 0.684 0.144 ;
      RECT 0.618 0.09 0.77 0.108 ;
      RECT 0.202 0.162 0.357 0.18 ;
      RECT 0.288 0.126 0.306 0.18 ;
      RECT 0.288 0.126 0.346 0.144 ;
      RECT 0.196 0.126 0.252 0.144 ;
      RECT 0.234 0.09 0.252 0.144 ;
      RECT 0.186 0.09 0.338 0.108 ;
  END
END CKINVDCx14_ASAP7_75t_L

MACRO CKINVDCx16_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx16_ASAP7_75t_L 0 0 ;
  SIZE 1.62 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.412 0.126 1.505 0.144 ;
        RECT 1.444 0.027 1.462 0.144 ;
        RECT 0.158 0.027 1.462 0.045 ;
        RECT 0.98 0.126 1.072 0.144 ;
        RECT 1.017 0.027 1.035 0.144 ;
        RECT 0.547 0.126 0.639 0.144 ;
        RECT 0.584 0.027 0.602 0.144 ;
        RECT 0.126 0.126 0.208 0.144 ;
        RECT 0.158 0.027 0.176 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.62 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.62 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.225 1.548 0.243 ;
        RECT 1.53 0.063 1.548 0.243 ;
        RECT 1.498 0.063 1.548 0.081 ;
        RECT 1.368 0.063 1.418 0.081 ;
        RECT 1.368 0.063 1.386 0.243 ;
        RECT 1.098 0.063 1.116 0.243 ;
        RECT 1.066 0.063 1.116 0.081 ;
        RECT 0.936 0.063 0.986 0.081 ;
        RECT 0.936 0.063 0.954 0.243 ;
        RECT 0.666 0.063 0.684 0.243 ;
        RECT 0.634 0.063 0.684 0.081 ;
        RECT 0.504 0.063 0.554 0.081 ;
        RECT 0.504 0.063 0.522 0.243 ;
        RECT 0.234 0.063 0.252 0.243 ;
        RECT 0.202 0.063 0.252 0.081 ;
        RECT 0.072 0.063 0.122 0.081 ;
        RECT 0.072 0.063 0.09 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.26 0.126 1.316 0.144 ;
      RECT 1.26 0.09 1.278 0.144 ;
      RECT 1.174 0.09 1.326 0.108 ;
      RECT 1.155 0.162 1.31 0.18 ;
      RECT 1.206 0.126 1.224 0.18 ;
      RECT 1.166 0.126 1.224 0.144 ;
      RECT 0.742 0.162 0.897 0.18 ;
      RECT 0.828 0.126 0.846 0.18 ;
      RECT 0.828 0.126 0.886 0.144 ;
      RECT 0.736 0.126 0.792 0.144 ;
      RECT 0.774 0.09 0.792 0.144 ;
      RECT 0.726 0.09 0.878 0.108 ;
      RECT 0.31 0.162 0.465 0.18 ;
      RECT 0.396 0.126 0.414 0.18 ;
      RECT 0.396 0.126 0.454 0.144 ;
      RECT 0.304 0.126 0.36 0.144 ;
      RECT 0.342 0.09 0.36 0.144 ;
      RECT 0.294 0.09 0.446 0.108 ;
  END
END CKINVDCx16_ASAP7_75t_L

MACRO CKINVDCx20_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx20_ASAP7_75t_L 0 0 ;
  SIZE 2.052 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.844 0.126 1.937 0.144 ;
        RECT 1.876 0.027 1.894 0.144 ;
        RECT 0.158 0.027 1.894 0.045 ;
        RECT 1.412 0.126 1.505 0.144 ;
        RECT 1.444 0.027 1.462 0.144 ;
        RECT 0.98 0.126 1.072 0.144 ;
        RECT 1.017 0.027 1.035 0.144 ;
        RECT 0.547 0.126 0.639 0.144 ;
        RECT 0.584 0.027 0.602 0.144 ;
        RECT 0.126 0.126 0.208 0.144 ;
        RECT 0.158 0.027 0.176 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.052 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.052 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.225 1.98 0.243 ;
        RECT 1.962 0.063 1.98 0.243 ;
        RECT 1.93 0.063 1.98 0.081 ;
        RECT 1.8 0.063 1.85 0.081 ;
        RECT 1.8 0.063 1.818 0.243 ;
        RECT 1.53 0.063 1.548 0.243 ;
        RECT 1.498 0.063 1.548 0.081 ;
        RECT 1.368 0.063 1.418 0.081 ;
        RECT 1.368 0.063 1.386 0.243 ;
        RECT 1.098 0.063 1.116 0.243 ;
        RECT 1.066 0.063 1.116 0.081 ;
        RECT 0.936 0.063 0.986 0.081 ;
        RECT 0.936 0.063 0.954 0.243 ;
        RECT 0.666 0.063 0.684 0.243 ;
        RECT 0.634 0.063 0.684 0.081 ;
        RECT 0.504 0.063 0.554 0.081 ;
        RECT 0.504 0.063 0.522 0.243 ;
        RECT 0.234 0.063 0.252 0.243 ;
        RECT 0.202 0.063 0.252 0.081 ;
        RECT 0.072 0.063 0.122 0.081 ;
        RECT 0.072 0.063 0.09 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.692 0.126 1.748 0.144 ;
      RECT 1.692 0.09 1.71 0.144 ;
      RECT 1.606 0.09 1.758 0.108 ;
      RECT 1.587 0.162 1.742 0.18 ;
      RECT 1.638 0.126 1.656 0.18 ;
      RECT 1.598 0.126 1.656 0.144 ;
      RECT 1.26 0.126 1.316 0.144 ;
      RECT 1.26 0.09 1.278 0.144 ;
      RECT 1.174 0.09 1.326 0.108 ;
      RECT 1.155 0.162 1.31 0.18 ;
      RECT 1.206 0.126 1.224 0.18 ;
      RECT 1.166 0.126 1.224 0.144 ;
      RECT 0.742 0.162 0.897 0.18 ;
      RECT 0.828 0.126 0.846 0.18 ;
      RECT 0.828 0.126 0.886 0.144 ;
      RECT 0.736 0.126 0.792 0.144 ;
      RECT 0.774 0.09 0.792 0.144 ;
      RECT 0.726 0.09 0.878 0.108 ;
      RECT 0.31 0.162 0.465 0.18 ;
      RECT 0.396 0.126 0.414 0.18 ;
      RECT 0.396 0.126 0.454 0.144 ;
      RECT 0.304 0.126 0.36 0.144 ;
      RECT 0.342 0.09 0.36 0.144 ;
      RECT 0.294 0.09 0.446 0.108 ;
  END
END CKINVDCx20_ASAP7_75t_L

MACRO CKINVDCx5p33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx5p33_ASAP7_75t_L 0 0 ;
  SIZE 1.188 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.088 0.126 1.138 0.144 ;
        RECT 1.12 0.027 1.138 0.144 ;
        RECT 0.05 0.027 1.138 0.045 ;
        RECT 0.764 0.126 0.814 0.144 ;
        RECT 0.796 0.027 0.814 0.144 ;
        RECT 0.374 0.126 0.424 0.144 ;
        RECT 0.374 0.027 0.392 0.144 ;
        RECT 0.05 0.126 0.1 0.144 ;
        RECT 0.05 0.027 0.068 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 1.094 0.243 ;
        RECT 1.044 0.063 1.094 0.081 ;
        RECT 1.044 0.063 1.062 0.243 ;
        RECT 0.72 0.063 0.77 0.081 ;
        RECT 0.72 0.063 0.738 0.243 ;
        RECT 0.45 0.063 0.468 0.243 ;
        RECT 0.418 0.063 0.468 0.081 ;
        RECT 0.126 0.063 0.144 0.243 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.936 0.126 0.992 0.144 ;
      RECT 0.936 0.09 0.954 0.144 ;
      RECT 0.85 0.09 1.002 0.108 ;
      RECT 0.831 0.162 0.986 0.18 ;
      RECT 0.882 0.126 0.9 0.18 ;
      RECT 0.842 0.126 0.9 0.144 ;
      RECT 0.526 0.162 0.681 0.18 ;
      RECT 0.612 0.126 0.63 0.18 ;
      RECT 0.612 0.126 0.67 0.144 ;
      RECT 0.52 0.126 0.576 0.144 ;
      RECT 0.558 0.09 0.576 0.144 ;
      RECT 0.51 0.09 0.662 0.108 ;
      RECT 0.202 0.162 0.357 0.18 ;
      RECT 0.288 0.126 0.306 0.18 ;
      RECT 0.288 0.126 0.346 0.144 ;
      RECT 0.196 0.126 0.252 0.144 ;
      RECT 0.234 0.09 0.252 0.144 ;
      RECT 0.186 0.09 0.338 0.108 ;
  END
END CKINVDCx5p33_ASAP7_75t_L

MACRO CKINVDCx6p67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx6p67_ASAP7_75t_L 0 0 ;
  SIZE 1.296 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.088 0.126 1.17 0.144 ;
        RECT 1.12 0.027 1.138 0.144 ;
        RECT 0.05 0.027 1.138 0.045 ;
        RECT 0.764 0.126 0.814 0.144 ;
        RECT 0.796 0.027 0.814 0.144 ;
        RECT 0.374 0.126 0.424 0.144 ;
        RECT 0.374 0.027 0.392 0.144 ;
        RECT 0.05 0.126 0.1 0.144 ;
        RECT 0.05 0.027 0.068 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.296 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.296 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 1.224 0.243 ;
        RECT 1.206 0.063 1.224 0.243 ;
        RECT 1.174 0.063 1.224 0.081 ;
        RECT 1.044 0.063 1.094 0.081 ;
        RECT 1.044 0.063 1.062 0.243 ;
        RECT 0.72 0.063 0.77 0.081 ;
        RECT 0.72 0.063 0.738 0.243 ;
        RECT 0.45 0.063 0.468 0.243 ;
        RECT 0.418 0.063 0.468 0.081 ;
        RECT 0.126 0.063 0.144 0.243 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.936 0.126 0.992 0.144 ;
      RECT 0.936 0.09 0.954 0.144 ;
      RECT 0.85 0.09 1.002 0.108 ;
      RECT 0.831 0.162 0.986 0.18 ;
      RECT 0.882 0.126 0.9 0.18 ;
      RECT 0.842 0.126 0.9 0.144 ;
      RECT 0.526 0.162 0.681 0.18 ;
      RECT 0.612 0.126 0.63 0.18 ;
      RECT 0.612 0.126 0.67 0.144 ;
      RECT 0.52 0.126 0.576 0.144 ;
      RECT 0.558 0.09 0.576 0.144 ;
      RECT 0.51 0.09 0.662 0.108 ;
      RECT 0.202 0.162 0.357 0.18 ;
      RECT 0.288 0.126 0.306 0.18 ;
      RECT 0.288 0.126 0.346 0.144 ;
      RECT 0.196 0.126 0.252 0.144 ;
      RECT 0.234 0.09 0.252 0.144 ;
      RECT 0.186 0.09 0.338 0.108 ;
  END
END CKINVDCx6p67_ASAP7_75t_L

MACRO CKINVDCx8_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx8_ASAP7_75t_L 0 0 ;
  SIZE 1.188 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.088 0.126 1.138 0.144 ;
        RECT 1.12 0.027 1.138 0.144 ;
        RECT 0.05 0.027 1.138 0.045 ;
        RECT 0.764 0.126 0.814 0.144 ;
        RECT 0.796 0.027 0.814 0.144 ;
        RECT 0.374 0.126 0.424 0.144 ;
        RECT 0.374 0.027 0.392 0.144 ;
        RECT 0.05 0.126 0.1 0.144 ;
        RECT 0.05 0.027 0.068 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 1.094 0.243 ;
        RECT 1.044 0.063 1.094 0.081 ;
        RECT 1.044 0.063 1.062 0.243 ;
        RECT 0.72 0.063 0.77 0.081 ;
        RECT 0.72 0.063 0.738 0.243 ;
        RECT 0.45 0.063 0.468 0.243 ;
        RECT 0.418 0.063 0.468 0.081 ;
        RECT 0.126 0.063 0.144 0.243 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.936 0.126 0.992 0.144 ;
      RECT 0.936 0.09 0.954 0.144 ;
      RECT 0.85 0.09 1.002 0.108 ;
      RECT 0.831 0.162 0.986 0.18 ;
      RECT 0.882 0.126 0.9 0.18 ;
      RECT 0.842 0.126 0.9 0.144 ;
      RECT 0.526 0.162 0.681 0.18 ;
      RECT 0.612 0.126 0.63 0.18 ;
      RECT 0.612 0.126 0.67 0.144 ;
      RECT 0.52 0.126 0.576 0.144 ;
      RECT 0.558 0.09 0.576 0.144 ;
      RECT 0.51 0.09 0.662 0.108 ;
      RECT 0.202 0.162 0.357 0.18 ;
      RECT 0.288 0.126 0.306 0.18 ;
      RECT 0.288 0.126 0.346 0.144 ;
      RECT 0.196 0.126 0.252 0.144 ;
      RECT 0.234 0.09 0.252 0.144 ;
      RECT 0.186 0.09 0.338 0.108 ;
  END
END CKINVDCx8_ASAP7_75t_L

MACRO CKINVDCx9p33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx9p33_ASAP7_75t_L 0 0 ;
  SIZE 1.512 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.304 0.126 1.397 0.144 ;
        RECT 1.336 0.027 1.354 0.144 ;
        RECT 0.05 0.027 1.354 0.045 ;
        RECT 0.872 0.126 0.964 0.144 ;
        RECT 0.909 0.027 0.927 0.144 ;
        RECT 0.439 0.126 0.531 0.144 ;
        RECT 0.476 0.027 0.494 0.144 ;
        RECT 0.05 0.126 0.1 0.144 ;
        RECT 0.05 0.027 0.068 0.144 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.512 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.512 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 1.44 0.243 ;
        RECT 1.422 0.063 1.44 0.243 ;
        RECT 1.39 0.063 1.44 0.081 ;
        RECT 1.26 0.063 1.31 0.081 ;
        RECT 1.26 0.063 1.278 0.243 ;
        RECT 0.99 0.063 1.008 0.243 ;
        RECT 0.958 0.063 1.008 0.081 ;
        RECT 0.828 0.063 0.878 0.081 ;
        RECT 0.828 0.063 0.846 0.243 ;
        RECT 0.558 0.063 0.576 0.243 ;
        RECT 0.526 0.063 0.576 0.081 ;
        RECT 0.396 0.063 0.446 0.081 ;
        RECT 0.396 0.063 0.414 0.243 ;
        RECT 0.126 0.063 0.144 0.243 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.152 0.126 1.208 0.144 ;
      RECT 1.152 0.09 1.17 0.144 ;
      RECT 1.066 0.09 1.218 0.108 ;
      RECT 1.047 0.162 1.202 0.18 ;
      RECT 1.098 0.126 1.116 0.18 ;
      RECT 1.058 0.126 1.116 0.144 ;
      RECT 0.634 0.162 0.789 0.18 ;
      RECT 0.72 0.126 0.738 0.18 ;
      RECT 0.72 0.126 0.778 0.144 ;
      RECT 0.628 0.126 0.684 0.144 ;
      RECT 0.666 0.09 0.684 0.144 ;
      RECT 0.618 0.09 0.77 0.108 ;
      RECT 0.202 0.162 0.357 0.18 ;
      RECT 0.288 0.126 0.306 0.18 ;
      RECT 0.288 0.126 0.346 0.144 ;
      RECT 0.196 0.126 0.252 0.144 ;
      RECT 0.234 0.09 0.252 0.144 ;
      RECT 0.186 0.09 0.338 0.108 ;
  END
END CKINVDCx9p33_ASAP7_75t_L

MACRO DECAPx10_ASAP7_75t_L
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx10_ASAP7_75t_L 0 0 ;
  SIZE 1.188 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.558 0.045 0.576 0.15 ;
      RECT 0.558 0.045 1.148 0.063 ;
      RECT 0.04 0.207 0.63 0.225 ;
      RECT 0.612 0.121 0.63 0.225 ;
  END
END DECAPx10_ASAP7_75t_L

MACRO DECAPx1_ASAP7_75t_L
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx1_ASAP7_75t_L 0 0 ;
  SIZE 0.216 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.216 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.094 0.207 0.144 0.225 ;
      RECT 0.126 0.121 0.144 0.225 ;
      RECT 0.072 0.045 0.09 0.15 ;
      RECT 0.072 0.045 0.122 0.063 ;
  END
END DECAPx1_ASAP7_75t_L

MACRO DECAPx2_ASAP7_75t_L
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx2_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.126 0.045 0.144 0.15 ;
      RECT 0.126 0.045 0.284 0.063 ;
      RECT 0.04 0.207 0.198 0.225 ;
      RECT 0.18 0.121 0.198 0.225 ;
  END
END DECAPx2_ASAP7_75t_L

MACRO DECAPx2b_ASAP7_75t_L
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx2b_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.094 0.162 0.249 0.18 ;
      RECT 0.18 0.126 0.198 0.18 ;
      RECT 0.18 0.126 0.238 0.144 ;
      RECT 0.088 0.126 0.144 0.144 ;
      RECT 0.126 0.09 0.144 0.144 ;
      RECT 0.078 0.09 0.23 0.108 ;
  END
END DECAPx2b_ASAP7_75t_L

MACRO DECAPx4_ASAP7_75t_L
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx4_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.234 0.045 0.252 0.15 ;
      RECT 0.234 0.045 0.5 0.063 ;
      RECT 0.04 0.207 0.306 0.225 ;
      RECT 0.288 0.121 0.306 0.225 ;
  END
END DECAPx4_ASAP7_75t_L

MACRO DECAPx6_ASAP7_75t_L
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx6_ASAP7_75t_L 0 0 ;
  SIZE 0.756 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.756 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.342 0.045 0.36 0.15 ;
      RECT 0.342 0.045 0.716 0.063 ;
      RECT 0.04 0.207 0.414 0.225 ;
      RECT 0.396 0.121 0.414 0.225 ;
  END
END DECAPx6_ASAP7_75t_L

MACRO DFFHQNx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx1_ASAP7_75t_L 0 0 ;
  SIZE 1.08 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.062 0.243 ;
        RECT 1.044 0.027 1.062 0.243 ;
        RECT 1.012 0.027 1.062 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.08 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.142 0.106 0.16 0.167 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.175 0.18 0.527 0.198 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END DFFHQNx1_ASAP7_75t_L

MACRO DFFHQNx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx2_ASAP7_75t_L 0 0 ;
  SIZE 1.134 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.216 1.117 0.234 ;
        RECT 1.099 0.036 1.117 0.234 ;
        RECT 1.012 0.036 1.117 0.054 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.134 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.134 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.142 0.106 0.16 0.167 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.175 0.18 0.527 0.198 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END DFFHQNx2_ASAP7_75t_L

MACRO DFFHQNx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx3_ASAP7_75t_L 0 0 ;
  SIZE 1.188 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.171 0.243 ;
        RECT 1.153 0.027 1.171 0.243 ;
        RECT 1.012 0.027 1.171 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.99 0.122 1.008 0.167 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.142 0.106 0.16 0.167 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.175 0.18 0.527 0.198 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END DFFHQNx3_ASAP7_75t_L

MACRO DFFHQx4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQx4_ASAP7_75t_L 0 0 ;
  SIZE 1.35 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.125 0.225 1.333 0.243 ;
        RECT 1.313 0.027 1.333 0.243 ;
        RECT 1.125 0.027 1.333 0.045 ;
        RECT 1.125 0.201 1.143 0.243 ;
        RECT 1.125 0.027 1.143 0.069 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.35 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.012 0.225 1.098 0.243 ;
      RECT 1.08 0.027 1.098 0.243 ;
      RECT 1.08 0.127 1.175 0.145 ;
      RECT 1.012 0.027 1.098 0.045 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.581 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.99 0.122 1.008 0.167 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.142 0.106 0.16 0.167 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.175 0.18 0.527 0.198 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END DFFHQx4_ASAP7_75t_L

MACRO DFFLQNx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQNx1_ASAP7_75t_L 0 0 ;
  SIZE 1.08 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.225 0.325 0.243 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.243 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.062 0.243 ;
        RECT 1.044 0.027 1.062 0.243 ;
        RECT 1.012 0.027 1.062 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.08 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.688 0.225 0.738 0.243 ;
      RECT 0.72 0.027 0.738 0.243 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.034 0.603 0.099 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.581 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.145 0.18 0.198 0.198 ;
      RECT 0.18 0.126 0.198 0.198 ;
      RECT 0.121 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.666 0.099 0.684 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.342 0.126 0.36 0.203 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.229 0.144 0.689 0.162 ;
      RECT 0.019 0.18 0.527 0.198 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.15 0.18 0.168 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END DFFLQNx1_ASAP7_75t_L

MACRO DFFLQNx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQNx2_ASAP7_75t_L 0 0 ;
  SIZE 1.134 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.115 0.243 ;
        RECT 1.097 0.027 1.115 0.243 ;
        RECT 1.012 0.027 1.115 0.045 ;
    END
  END QN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.225 0.325 0.243 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.243 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.134 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.134 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.688 0.225 0.738 0.243 ;
      RECT 0.72 0.027 0.738 0.243 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.034 0.603 0.099 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.581 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.145 0.18 0.198 0.198 ;
      RECT 0.18 0.126 0.198 0.198 ;
      RECT 0.121 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.666 0.099 0.684 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.342 0.126 0.36 0.203 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.229 0.144 0.689 0.162 ;
      RECT 0.019 0.18 0.527 0.198 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.15 0.18 0.168 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END DFFLQNx2_ASAP7_75t_L

MACRO DFFLQNx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQNx3_ASAP7_75t_L 0 0 ;
  SIZE 1.188 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.225 0.325 0.243 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.243 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.171 0.243 ;
        RECT 1.153 0.027 1.171 0.243 ;
        RECT 1.011 0.027 1.171 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.688 0.225 0.738 0.243 ;
      RECT 0.72 0.027 0.738 0.243 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.034 0.603 0.099 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.581 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.145 0.18 0.198 0.198 ;
      RECT 0.18 0.126 0.198 0.198 ;
      RECT 0.121 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.666 0.099 0.684 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.342 0.126 0.36 0.203 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.229 0.144 0.689 0.162 ;
      RECT 0.019 0.18 0.527 0.198 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.15 0.18 0.168 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END DFFLQNx3_ASAP7_75t_L

MACRO DFFLQx4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQx4_ASAP7_75t_L 0 0 ;
  SIZE 1.35 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.225 0.325 0.243 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.243 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.125 0.225 1.333 0.243 ;
        RECT 1.313 0.027 1.333 0.243 ;
        RECT 1.125 0.027 1.333 0.045 ;
        RECT 1.125 0.201 1.143 0.243 ;
        RECT 1.125 0.027 1.143 0.069 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.35 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.012 0.225 1.098 0.243 ;
      RECT 1.08 0.027 1.098 0.243 ;
      RECT 1.08 0.127 1.175 0.145 ;
      RECT 1.012 0.027 1.098 0.045 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.688 0.225 0.738 0.243 ;
      RECT 0.72 0.027 0.738 0.243 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.034 0.603 0.099 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.581 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.145 0.18 0.198 0.198 ;
      RECT 0.18 0.126 0.198 0.198 ;
      RECT 0.121 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.99 0.122 1.008 0.167 ;
      RECT 0.666 0.099 0.684 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.342 0.126 0.36 0.203 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.229 0.144 0.689 0.162 ;
      RECT 0.019 0.18 0.527 0.198 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.15 0.18 0.168 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END DFFLQx4_ASAP7_75t_L

MACRO DHLx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx1_ASAP7_75t_L 0 0 ;
  SIZE 0.81 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.153 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.117 ;
        RECT 0.099 0.034 0.117 0.117 ;
        RECT 0.072 0.153 0.117 0.189 ;
        RECT 0.072 0.081 0.09 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.236 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.742 0.225 0.792 0.243 ;
        RECT 0.774 0.027 0.792 0.243 ;
        RECT 0.742 0.027 0.792 0.045 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.81 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.58 0.225 0.63 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.504 0.027 0.522 0.096 ;
      RECT 0.504 0.027 0.63 0.045 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.121 0.581 0.139 ;
      RECT 0.414 0.027 0.468 0.045 ;
      RECT 0.342 0.189 0.379 0.207 ;
      RECT 0.342 0.106 0.36 0.207 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.148 0.18 0.198 0.198 ;
      RECT 0.18 0.126 0.198 0.198 ;
      RECT 0.138 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.72 0.122 0.738 0.167 ;
      RECT 0.504 0.164 0.522 0.207 ;
      RECT 0.396 0.106 0.414 0.171 ;
    LAYER M2 ;
      RECT 0.45 0.144 0.743 0.162 ;
      RECT 0.019 0.18 0.527 0.198 ;
      RECT 0.229 0.144 0.414 0.162 ;
    LAYER V1 ;
      RECT 0.72 0.144 0.738 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.153 0.18 0.171 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END DHLx1_ASAP7_75t_L

MACRO DHLx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx2_ASAP7_75t_L 0 0 ;
  SIZE 0.864 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.153 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.117 ;
        RECT 0.099 0.034 0.117 0.117 ;
        RECT 0.072 0.153 0.117 0.189 ;
        RECT 0.072 0.081 0.09 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.236 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.216 0.85 0.234 ;
        RECT 0.832 0.036 0.85 0.234 ;
        RECT 0.742 0.036 0.85 0.054 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.864 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.58 0.225 0.63 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.504 0.027 0.522 0.096 ;
      RECT 0.504 0.027 0.63 0.045 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.121 0.581 0.139 ;
      RECT 0.414 0.027 0.468 0.045 ;
      RECT 0.342 0.189 0.379 0.207 ;
      RECT 0.342 0.106 0.36 0.207 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.148 0.18 0.198 0.198 ;
      RECT 0.18 0.126 0.198 0.198 ;
      RECT 0.138 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.774 0.09 0.792 0.167 ;
      RECT 0.72 0.09 0.738 0.167 ;
      RECT 0.504 0.164 0.522 0.207 ;
      RECT 0.396 0.106 0.414 0.171 ;
    LAYER M2 ;
      RECT 0.45 0.144 0.797 0.162 ;
      RECT 0.019 0.18 0.527 0.198 ;
      RECT 0.229 0.144 0.414 0.162 ;
    LAYER V1 ;
      RECT 0.774 0.144 0.792 0.162 ;
      RECT 0.72 0.144 0.738 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.153 0.18 0.171 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END DHLx2_ASAP7_75t_L

MACRO DHLx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx3_ASAP7_75t_L 0 0 ;
  SIZE 0.918 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.153 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.117 ;
        RECT 0.099 0.034 0.117 0.117 ;
        RECT 0.072 0.153 0.117 0.189 ;
        RECT 0.072 0.081 0.09 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.236 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.688 0.225 0.9 0.243 ;
        RECT 0.882 0.027 0.9 0.243 ;
        RECT 0.688 0.027 0.9 0.045 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.918 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.918 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.58 0.225 0.63 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.504 0.027 0.522 0.096 ;
      RECT 0.504 0.027 0.63 0.045 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.121 0.581 0.139 ;
      RECT 0.414 0.027 0.468 0.045 ;
      RECT 0.342 0.189 0.379 0.207 ;
      RECT 0.342 0.106 0.36 0.207 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.148 0.18 0.198 0.198 ;
      RECT 0.18 0.126 0.198 0.198 ;
      RECT 0.138 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.828 0.09 0.846 0.167 ;
      RECT 0.774 0.09 0.792 0.167 ;
      RECT 0.72 0.09 0.738 0.167 ;
      RECT 0.504 0.164 0.522 0.207 ;
      RECT 0.396 0.106 0.414 0.171 ;
    LAYER M2 ;
      RECT 0.45 0.144 0.851 0.162 ;
      RECT 0.019 0.18 0.527 0.198 ;
      RECT 0.229 0.144 0.414 0.162 ;
    LAYER V1 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.774 0.144 0.792 0.162 ;
      RECT 0.72 0.144 0.738 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.153 0.18 0.171 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END DHLx3_ASAP7_75t_L

MACRO DLLx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLLx1_ASAP7_75t_L 0 0 ;
  SIZE 0.81 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.153 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.117 ;
        RECT 0.099 0.034 0.117 0.117 ;
        RECT 0.072 0.153 0.117 0.189 ;
        RECT 0.072 0.081 0.09 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.225 0.325 0.243 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.243 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.742 0.225 0.792 0.243 ;
        RECT 0.774 0.027 0.792 0.243 ;
        RECT 0.735 0.027 0.792 0.045 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.81 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.58 0.225 0.63 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.504 0.027 0.522 0.097 ;
      RECT 0.504 0.027 0.63 0.045 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.58 0.14 ;
      RECT 0.414 0.027 0.468 0.045 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.148 0.189 0.198 0.207 ;
      RECT 0.18 0.126 0.198 0.207 ;
      RECT 0.138 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.72 0.106 0.738 0.2 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.2 ;
      RECT 0.342 0.106 0.36 0.203 ;
    LAYER M2 ;
      RECT 0.45 0.144 0.743 0.162 ;
      RECT 0.229 0.18 0.527 0.198 ;
      RECT 0.019 0.144 0.414 0.162 ;
    LAYER V1 ;
      RECT 0.72 0.144 0.738 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.18 0.252 0.198 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END DLLx1_ASAP7_75t_L

MACRO DLLx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLLx2_ASAP7_75t_L 0 0 ;
  SIZE 0.864 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.153 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.117 ;
        RECT 0.099 0.034 0.117 0.117 ;
        RECT 0.072 0.153 0.117 0.189 ;
        RECT 0.072 0.081 0.09 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.225 0.325 0.243 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.243 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.688 0.225 0.847 0.243 ;
        RECT 0.829 0.027 0.847 0.243 ;
        RECT 0.688 0.027 0.847 0.045 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.864 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.58 0.225 0.63 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.504 0.027 0.522 0.097 ;
      RECT 0.504 0.027 0.63 0.045 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.58 0.14 ;
      RECT 0.414 0.027 0.468 0.045 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.148 0.189 0.198 0.207 ;
      RECT 0.18 0.126 0.198 0.207 ;
      RECT 0.138 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.774 0.09 0.792 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.2 ;
      RECT 0.342 0.106 0.36 0.203 ;
    LAYER M2 ;
      RECT 0.45 0.144 0.8 0.162 ;
      RECT 0.229 0.18 0.527 0.198 ;
      RECT 0.019 0.144 0.414 0.162 ;
    LAYER V1 ;
      RECT 0.774 0.144 0.792 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.18 0.252 0.198 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END DLLx2_ASAP7_75t_L

MACRO DLLx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLLx3_ASAP7_75t_L 0 0 ;
  SIZE 0.918 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.153 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.117 ;
        RECT 0.099 0.034 0.117 0.117 ;
        RECT 0.072 0.153 0.117 0.189 ;
        RECT 0.072 0.081 0.09 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.225 0.325 0.243 ;
        RECT 0.288 0.027 0.325 0.045 ;
        RECT 0.288 0.027 0.306 0.243 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.742 0.216 0.901 0.234 ;
        RECT 0.882 0.036 0.901 0.234 ;
        RECT 0.742 0.036 0.901 0.054 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.918 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.918 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.58 0.225 0.63 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.504 0.027 0.522 0.097 ;
      RECT 0.504 0.027 0.63 0.045 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.58 0.14 ;
      RECT 0.414 0.027 0.468 0.045 ;
      RECT 0.148 0.225 0.252 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.148 0.189 0.198 0.207 ;
      RECT 0.18 0.126 0.198 0.207 ;
      RECT 0.138 0.126 0.198 0.144 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.774 0.09 0.792 0.167 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.396 0.106 0.414 0.2 ;
      RECT 0.342 0.106 0.36 0.203 ;
    LAYER M2 ;
      RECT 0.45 0.144 0.8 0.162 ;
      RECT 0.229 0.18 0.527 0.198 ;
      RECT 0.019 0.144 0.414 0.162 ;
    LAYER V1 ;
      RECT 0.774 0.144 0.792 0.162 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.342 0.18 0.36 0.198 ;
      RECT 0.234 0.18 0.252 0.198 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END DLLx3_ASAP7_75t_L

MACRO FAx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FAx1_ASAP7_75t_L 0 0 ;
  SIZE 0.756 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.324 0.225 0.495 0.243 ;
        RECT 0.477 0.184 0.495 0.243 ;
        RECT 0.477 0.027 0.495 0.068 ;
        RECT 0.324 0.027 0.495 0.045 ;
        RECT 0.324 0.027 0.342 0.243 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.756 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.059 0.18 0.627 0.198 ;
      LAYER M1 ;
        RECT 0.599 0.18 0.63 0.198 ;
        RECT 0.612 0.121 0.63 0.198 ;
        RECT 0.383 0.18 0.414 0.198 ;
        RECT 0.396 0.121 0.414 0.198 ;
        RECT 0.059 0.18 0.09 0.198 ;
        RECT 0.072 0.121 0.09 0.198 ;
      LAYER V1 ;
        RECT 0.064 0.18 0.082 0.198 ;
        RECT 0.388 0.18 0.406 0.198 ;
        RECT 0.604 0.18 0.622 0.198 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.167 0.144 0.689 0.162 ;
      LAYER M1 ;
        RECT 0.666 0.121 0.684 0.167 ;
        RECT 0.288 0.121 0.306 0.167 ;
        RECT 0.167 0.144 0.198 0.162 ;
        RECT 0.18 0.121 0.198 0.162 ;
      LAYER V1 ;
        RECT 0.172 0.144 0.19 0.162 ;
        RECT 0.288 0.144 0.306 0.162 ;
        RECT 0.666 0.144 0.684 0.162 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.229 0.108 0.587 0.126 ;
      LAYER M1 ;
        RECT 0.558 0.108 0.587 0.126 ;
        RECT 0.558 0.108 0.576 0.149 ;
        RECT 0.45 0.103 0.468 0.149 ;
        RECT 0.226 0.108 0.263 0.126 ;
        RECT 0.234 0.108 0.252 0.149 ;
      LAYER V1 ;
        RECT 0.234 0.108 0.252 0.126 ;
        RECT 0.45 0.108 0.468 0.126 ;
        RECT 0.564 0.108 0.582 0.126 ;
    END
  END CI
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.128 0.072 0.543 0.09 ;
      LAYER M1 ;
        RECT 0.515 0.072 0.543 0.09 ;
        RECT 0.504 0.09 0.533 0.108 ;
        RECT 0.504 0.09 0.522 0.149 ;
        RECT 0.124 0.072 0.282 0.09 ;
        RECT 0.124 0.189 0.23 0.207 ;
        RECT 0.124 0.072 0.142 0.207 ;
      LAYER V1 ;
        RECT 0.133 0.072 0.151 0.09 ;
        RECT 0.52 0.072 0.538 0.09 ;
    END
  END CON
  OBS
    LAYER M1 ;
      RECT 0.526 0.027 0.662 0.045 ;
      RECT 0.526 0.225 0.662 0.243 ;
      RECT 0.04 0.027 0.284 0.045 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END FAx1_ASAP7_75t_L

MACRO FILLER_ASAP7_75t_L
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLER_ASAP7_75t_L 0 0 ;
  SIZE 0.108 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.108 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.108 0.009 ;
    END
  END VSS
END FILLER_ASAP7_75t_L

MACRO FILLERxp5_ASAP7_75t_L
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLERxp5_ASAP7_75t_L 0 0 ;
  SIZE 0.054 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.054 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.054 0.009 ;
    END
  END VSS
END FILLERxp5_ASAP7_75t_L

MACRO HAxp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HAxp5_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.063 0.36 0.15 ;
        RECT 0.207 0.063 0.36 0.081 ;
        RECT 0.207 0.027 0.225 0.081 ;
        RECT 0.018 0.027 0.225 0.045 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.027 0.036 0.236 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.106 0.063 0.144 0.081 ;
    END
  END B
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.162 0.189 0.414 0.207 ;
        RECT 0.396 0.121 0.414 0.207 ;
        RECT 0.094 0.225 0.18 0.243 ;
        RECT 0.162 0.075 0.18 0.243 ;
    END
  END CON
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.423 0.027 0.468 0.045 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.256 0.027 0.387 0.045 ;
  END
END HAxp5_ASAP7_75t_L

MACRO HB1xp67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB1xp67_ASAP7_75t_L 0 0 ;
  SIZE 0.216 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.207 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.216 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.225 0.198 0.243 ;
        RECT 0.18 0.027 0.198 0.243 ;
        RECT 0.148 0.027 0.198 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.117 0.243 ;
      RECT 0.099 0.153 0.117 0.243 ;
      RECT 0.099 0.153 0.144 0.171 ;
      RECT 0.126 0.099 0.144 0.171 ;
      RECT 0.099 0.099 0.144 0.117 ;
      RECT 0.099 0.027 0.117 0.117 ;
      RECT 0.04 0.027 0.117 0.045 ;
  END
END HB1xp67_ASAP7_75t_L

MACRO HB2xp67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB2xp67_ASAP7_75t_L 0 0 ;
  SIZE 0.27 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.207 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.27 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.225 0.252 0.243 ;
        RECT 0.234 0.027 0.252 0.243 ;
        RECT 0.202 0.027 0.252 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.144 0.243 ;
      RECT 0.126 0.027 0.144 0.243 ;
      RECT 0.126 0.126 0.203 0.144 ;
      RECT 0.04 0.027 0.144 0.045 ;
  END
END HB2xp67_ASAP7_75t_L

MACRO HB3xp67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB3xp67_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.207 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.225 0.306 0.243 ;
        RECT 0.288 0.027 0.306 0.243 ;
        RECT 0.256 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.18 0.126 0.257 0.144 ;
      RECT 0.04 0.027 0.198 0.045 ;
  END
END HB3xp67_ASAP7_75t_L

MACRO HB4xp67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB4xp67_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.081 0.055 0.099 ;
        RECT 0.018 0.081 0.036 0.207 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.225 0.36 0.243 ;
        RECT 0.342 0.027 0.36 0.243 ;
        RECT 0.31 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.18 0.126 0.311 0.144 ;
      RECT 0.04 0.027 0.198 0.045 ;
  END
END HB4xp67_ASAP7_75t_L

MACRO ICGx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx1_ASAP7_75t_L 0 0 ;
  SIZE 0.972 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.199 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.899 0.225 0.954 0.243 ;
        RECT 0.936 0.027 0.954 0.243 ;
        RECT 0.879 0.027 0.954 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.199 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.972 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.972 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.229 0.144 0.635 0.162 ;
      LAYER M1 ;
        RECT 0.612 0.178 0.765 0.196 ;
        RECT 0.747 0.142 0.765 0.196 ;
        RECT 0.612 0.116 0.63 0.196 ;
        RECT 0.396 0.144 0.447 0.162 ;
        RECT 0.396 0.12 0.414 0.162 ;
        RECT 0.234 0.119 0.252 0.184 ;
      LAYER V1 ;
        RECT 0.234 0.144 0.252 0.162 ;
        RECT 0.414 0.144 0.432 0.162 ;
        RECT 0.612 0.144 0.63 0.162 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.688 0.222 0.846 0.24 ;
      RECT 0.828 0.188 0.846 0.24 ;
      RECT 0.828 0.188 0.9 0.206 ;
      RECT 0.882 0.063 0.9 0.206 ;
      RECT 0.742 0.063 0.9 0.081 ;
      RECT 0.256 0.223 0.367 0.241 ;
      RECT 0.349 0.027 0.367 0.241 ;
      RECT 0.349 0.181 0.473 0.199 ;
      RECT 0.828 0.099 0.846 0.147 ;
      RECT 0.666 0.027 0.684 0.147 ;
      RECT 0.666 0.099 0.846 0.117 ;
      RECT 0.31 0.027 0.684 0.045 ;
      RECT 0.559 0.223 0.609 0.241 ;
      RECT 0.559 0.077 0.577 0.241 ;
      RECT 0.559 0.077 0.609 0.095 ;
      RECT 0.468 0.224 0.522 0.242 ;
      RECT 0.503 0.073 0.522 0.242 ;
      RECT 0.392 0.073 0.522 0.091 ;
      RECT 0.288 0.18 0.324 0.198 ;
      RECT 0.288 0.072 0.306 0.198 ;
      RECT 0.037 0.224 0.198 0.242 ;
      RECT 0.18 0.027 0.198 0.242 ;
      RECT 0.089 0.027 0.198 0.045 ;
    LAYER M2 ;
      RECT 0.296 0.18 0.582 0.198 ;
    LAYER V1 ;
      RECT 0.559 0.18 0.577 0.198 ;
      RECT 0.301 0.18 0.319 0.198 ;
  END
END ICGx1_ASAP7_75t_L

MACRO ICGx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx2_ASAP7_75t_L 0 0 ;
  SIZE 1.026 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.199 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.899 0.225 1.008 0.243 ;
        RECT 0.99 0.027 1.008 0.243 ;
        RECT 0.879 0.027 1.008 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.199 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.026 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.026 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.229 0.144 0.635 0.162 ;
      LAYER M1 ;
        RECT 0.612 0.178 0.765 0.196 ;
        RECT 0.747 0.142 0.765 0.196 ;
        RECT 0.612 0.116 0.63 0.196 ;
        RECT 0.396 0.144 0.447 0.162 ;
        RECT 0.396 0.12 0.414 0.162 ;
        RECT 0.234 0.119 0.252 0.184 ;
      LAYER V1 ;
        RECT 0.234 0.144 0.252 0.162 ;
        RECT 0.414 0.144 0.432 0.162 ;
        RECT 0.612 0.144 0.63 0.162 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.688 0.222 0.846 0.24 ;
      RECT 0.828 0.188 0.846 0.24 ;
      RECT 0.828 0.188 0.9 0.206 ;
      RECT 0.882 0.063 0.9 0.206 ;
      RECT 0.742 0.063 0.9 0.081 ;
      RECT 0.256 0.223 0.367 0.241 ;
      RECT 0.349 0.027 0.367 0.241 ;
      RECT 0.349 0.181 0.473 0.199 ;
      RECT 0.828 0.099 0.846 0.147 ;
      RECT 0.666 0.027 0.684 0.147 ;
      RECT 0.666 0.099 0.846 0.117 ;
      RECT 0.31 0.027 0.684 0.045 ;
      RECT 0.559 0.223 0.609 0.241 ;
      RECT 0.559 0.077 0.577 0.241 ;
      RECT 0.559 0.077 0.609 0.095 ;
      RECT 0.468 0.224 0.522 0.242 ;
      RECT 0.503 0.073 0.522 0.242 ;
      RECT 0.392 0.073 0.522 0.091 ;
      RECT 0.288 0.18 0.324 0.198 ;
      RECT 0.288 0.072 0.306 0.198 ;
      RECT 0.257 0.072 0.306 0.09 ;
      RECT 0.037 0.224 0.198 0.242 ;
      RECT 0.18 0.027 0.198 0.242 ;
      RECT 0.089 0.027 0.198 0.045 ;
    LAYER M2 ;
      RECT 0.296 0.18 0.582 0.198 ;
    LAYER V1 ;
      RECT 0.559 0.18 0.577 0.198 ;
      RECT 0.301 0.18 0.319 0.198 ;
  END
END ICGx2_ASAP7_75t_L

MACRO ICGx2p67DC_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx2p67DC_ASAP7_75t_L 0 0 ;
  SIZE 2.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.466 0.225 2.521 0.243 ;
        RECT 2.503 0.027 2.521 0.243 ;
        RECT 2.446 0.027 2.521 0.045 ;
        RECT 1.926 0.225 1.981 0.243 ;
        RECT 1.963 0.027 1.981 0.243 ;
        RECT 1.906 0.027 1.981 0.045 ;
        RECT 0.613 0.027 0.688 0.045 ;
        RECT 0.613 0.225 0.668 0.243 ;
        RECT 0.613 0.027 0.631 0.243 ;
        RECT 0.073 0.027 0.148 0.045 ;
        RECT 0.073 0.225 0.128 0.243 ;
        RECT 0.073 0.027 0.091 0.243 ;
      LAYER M2 ;
        RECT 0.062 0.036 2.532 0.054 ;
      LAYER V1 ;
        RECT 0.073 0.036 0.091 0.054 ;
        RECT 0.613 0.036 0.631 0.054 ;
        RECT 1.963 0.036 1.981 0.054 ;
        RECT 2.503 0.036 2.521 0.054 ;
    END
  END GCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.594 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 2.282 0.171 2.351 0.189 ;
        RECT 2.333 0.135 2.351 0.189 ;
        RECT 2.293 0.135 2.351 0.153 ;
        RECT 1.639 0.178 1.792 0.196 ;
        RECT 1.774 0.142 1.792 0.196 ;
        RECT 1.639 0.116 1.657 0.196 ;
        RECT 1.423 0.144 1.474 0.162 ;
        RECT 1.423 0.12 1.441 0.162 ;
        RECT 1.261 0.119 1.279 0.184 ;
        RECT 0.802 0.178 0.955 0.196 ;
        RECT 0.937 0.116 0.955 0.196 ;
        RECT 0.802 0.142 0.82 0.196 ;
        RECT 0.249 0.171 0.318 0.189 ;
        RECT 0.249 0.135 0.307 0.153 ;
        RECT 0.249 0.135 0.267 0.189 ;
      LAYER M2 ;
        RECT 0.236 0.144 2.359 0.162 ;
      LAYER V1 ;
        RECT 0.249 0.144 0.267 0.162 ;
        RECT 0.937 0.144 0.955 0.162 ;
        RECT 1.261 0.144 1.279 0.162 ;
        RECT 1.441 0.144 1.459 0.162 ;
        RECT 1.639 0.144 1.657 0.162 ;
        RECT 2.333 0.144 2.351 0.162 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.077 0.172 1.117 0.199 ;
        RECT 1.099 0.07 1.117 0.199 ;
        RECT 1.033 0.222 1.096 0.241 ;
        RECT 1.077 0.172 1.096 0.241 ;
      LAYER M2 ;
        RECT 0.983 0.216 1.238 0.234 ;
      LAYER V1 ;
        RECT 1.077 0.216 1.096 0.234 ;
    END
  END ENA
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.153 0.07 1.171 0.199 ;
      LAYER M2 ;
        RECT 0.983 0.072 1.238 0.09 ;
      LAYER V1 ;
        RECT 1.153 0.072 1.171 0.09 ;
    END
  END SE
  OBS
    LAYER M1 ;
      RECT 2.255 0.222 2.413 0.24 ;
      RECT 2.395 0.188 2.413 0.24 ;
      RECT 2.395 0.188 2.467 0.206 ;
      RECT 2.449 0.063 2.467 0.206 ;
      RECT 2.309 0.063 2.467 0.081 ;
      RECT 2.395 0.099 2.413 0.147 ;
      RECT 2.233 0.099 2.251 0.147 ;
      RECT 2.233 0.099 2.413 0.117 ;
      RECT 2.125 0.126 2.181 0.144 ;
      RECT 2.125 0.09 2.143 0.144 ;
      RECT 2.039 0.09 2.191 0.108 ;
      RECT 2.02 0.162 2.175 0.18 ;
      RECT 2.071 0.126 2.089 0.18 ;
      RECT 2.031 0.126 2.089 0.144 ;
      RECT 1.715 0.222 1.873 0.24 ;
      RECT 1.855 0.188 1.873 0.24 ;
      RECT 1.855 0.188 1.927 0.206 ;
      RECT 1.909 0.063 1.927 0.206 ;
      RECT 1.769 0.063 1.927 0.081 ;
      RECT 1.283 0.223 1.394 0.241 ;
      RECT 1.376 0.027 1.394 0.241 ;
      RECT 1.376 0.181 1.5 0.199 ;
      RECT 1.855 0.099 1.873 0.147 ;
      RECT 1.693 0.027 1.711 0.147 ;
      RECT 1.693 0.099 1.873 0.117 ;
      RECT 1.337 0.027 1.711 0.045 ;
      RECT 1.586 0.223 1.636 0.241 ;
      RECT 1.586 0.077 1.604 0.241 ;
      RECT 1.586 0.077 1.636 0.095 ;
      RECT 1.495 0.224 1.549 0.242 ;
      RECT 1.53 0.073 1.549 0.242 ;
      RECT 1.419 0.073 1.549 0.091 ;
      RECT 1.315 0.18 1.351 0.198 ;
      RECT 1.315 0.072 1.333 0.198 ;
      RECT 1.284 0.072 1.333 0.09 ;
      RECT 1.121 0.224 1.225 0.242 ;
      RECT 1.207 0.027 1.225 0.242 ;
      RECT 1.116 0.027 1.225 0.045 ;
      RECT 0.958 0.223 1.008 0.241 ;
      RECT 0.99 0.077 1.008 0.241 ;
      RECT 0.958 0.077 1.008 0.095 ;
      RECT 0.883 0.099 0.901 0.147 ;
      RECT 0.721 0.099 0.739 0.147 ;
      RECT 0.721 0.099 0.901 0.117 ;
      RECT 0.721 0.222 0.879 0.24 ;
      RECT 0.721 0.188 0.739 0.24 ;
      RECT 0.667 0.188 0.739 0.206 ;
      RECT 0.667 0.063 0.685 0.206 ;
      RECT 0.667 0.063 0.825 0.081 ;
      RECT 0.419 0.162 0.574 0.18 ;
      RECT 0.505 0.126 0.523 0.18 ;
      RECT 0.505 0.126 0.563 0.144 ;
      RECT 0.413 0.126 0.469 0.144 ;
      RECT 0.451 0.09 0.469 0.144 ;
      RECT 0.403 0.09 0.555 0.108 ;
      RECT 0.343 0.099 0.361 0.147 ;
      RECT 0.181 0.099 0.199 0.147 ;
      RECT 0.181 0.099 0.361 0.117 ;
      RECT 0.181 0.222 0.339 0.24 ;
      RECT 0.181 0.188 0.199 0.24 ;
      RECT 0.127 0.188 0.199 0.206 ;
      RECT 0.127 0.063 0.145 0.206 ;
      RECT 0.127 0.063 0.285 0.081 ;
    LAYER M2 ;
      RECT 0.337 0.108 2.257 0.126 ;
      RECT 0.983 0.18 1.609 0.198 ;
    LAYER V1 ;
      RECT 2.233 0.108 2.251 0.126 ;
      RECT 1.693 0.108 1.711 0.126 ;
      RECT 1.586 0.18 1.604 0.198 ;
      RECT 1.328 0.18 1.346 0.198 ;
      RECT 0.99 0.18 1.008 0.198 ;
      RECT 0.883 0.108 0.901 0.126 ;
      RECT 0.343 0.108 0.361 0.126 ;
  END
END ICGx2p67DC_ASAP7_75t_L

MACRO ICGx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx3_ASAP7_75t_L 0 0 ;
  SIZE 1.08 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.199 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.899 0.225 1.062 0.243 ;
        RECT 1.044 0.027 1.062 0.243 ;
        RECT 0.879 0.027 1.062 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.199 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.08 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.229 0.144 0.635 0.162 ;
      LAYER M1 ;
        RECT 0.612 0.178 0.765 0.196 ;
        RECT 0.747 0.142 0.765 0.196 ;
        RECT 0.612 0.116 0.63 0.196 ;
        RECT 0.396 0.144 0.447 0.162 ;
        RECT 0.396 0.12 0.414 0.162 ;
        RECT 0.234 0.119 0.252 0.184 ;
      LAYER V1 ;
        RECT 0.234 0.144 0.252 0.162 ;
        RECT 0.414 0.144 0.432 0.162 ;
        RECT 0.612 0.144 0.63 0.162 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.688 0.222 0.846 0.24 ;
      RECT 0.828 0.188 0.846 0.24 ;
      RECT 0.828 0.188 0.9 0.206 ;
      RECT 0.882 0.063 0.9 0.206 ;
      RECT 0.742 0.063 0.9 0.081 ;
      RECT 0.256 0.223 0.367 0.241 ;
      RECT 0.349 0.027 0.367 0.241 ;
      RECT 0.349 0.181 0.473 0.199 ;
      RECT 0.828 0.099 0.846 0.147 ;
      RECT 0.666 0.027 0.684 0.147 ;
      RECT 0.666 0.099 0.846 0.117 ;
      RECT 0.31 0.027 0.684 0.045 ;
      RECT 0.559 0.223 0.609 0.241 ;
      RECT 0.559 0.077 0.577 0.241 ;
      RECT 0.559 0.077 0.609 0.095 ;
      RECT 0.468 0.224 0.522 0.242 ;
      RECT 0.503 0.073 0.522 0.242 ;
      RECT 0.392 0.073 0.522 0.091 ;
      RECT 0.288 0.18 0.324 0.198 ;
      RECT 0.288 0.072 0.306 0.198 ;
      RECT 0.257 0.072 0.306 0.09 ;
      RECT 0.037 0.224 0.198 0.242 ;
      RECT 0.18 0.027 0.198 0.242 ;
      RECT 0.089 0.027 0.198 0.045 ;
    LAYER M2 ;
      RECT 0.296 0.18 0.582 0.198 ;
    LAYER V1 ;
      RECT 0.559 0.18 0.577 0.198 ;
      RECT 0.301 0.18 0.319 0.198 ;
  END
END ICGx3_ASAP7_75t_L

MACRO ICGx4DC_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx4DC_ASAP7_75t_L 0 0 ;
  SIZE 2.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.466 0.225 2.521 0.243 ;
        RECT 2.503 0.027 2.521 0.243 ;
        RECT 2.446 0.027 2.521 0.045 ;
        RECT 1.926 0.225 1.981 0.243 ;
        RECT 1.963 0.027 1.981 0.243 ;
        RECT 1.906 0.027 1.981 0.045 ;
        RECT 0.613 0.027 0.688 0.045 ;
        RECT 0.613 0.225 0.668 0.243 ;
        RECT 0.613 0.027 0.631 0.243 ;
        RECT 0.073 0.027 0.148 0.045 ;
        RECT 0.073 0.225 0.128 0.243 ;
        RECT 0.073 0.027 0.091 0.243 ;
      LAYER M2 ;
        RECT 0.062 0.036 2.532 0.054 ;
      LAYER V1 ;
        RECT 0.073 0.036 0.091 0.054 ;
        RECT 0.613 0.036 0.631 0.054 ;
        RECT 1.963 0.036 1.981 0.054 ;
        RECT 2.503 0.036 2.521 0.054 ;
    END
  END GCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.594 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 2.282 0.171 2.351 0.189 ;
        RECT 2.333 0.135 2.351 0.189 ;
        RECT 2.293 0.135 2.351 0.153 ;
        RECT 1.639 0.178 1.792 0.196 ;
        RECT 1.774 0.142 1.792 0.196 ;
        RECT 1.639 0.116 1.657 0.196 ;
        RECT 1.423 0.144 1.474 0.162 ;
        RECT 1.423 0.12 1.441 0.162 ;
        RECT 1.261 0.119 1.279 0.184 ;
        RECT 0.802 0.178 0.955 0.196 ;
        RECT 0.937 0.116 0.955 0.196 ;
        RECT 0.802 0.142 0.82 0.196 ;
        RECT 0.249 0.171 0.318 0.189 ;
        RECT 0.249 0.135 0.307 0.153 ;
        RECT 0.249 0.135 0.267 0.189 ;
      LAYER M2 ;
        RECT 0.236 0.144 2.359 0.162 ;
      LAYER V1 ;
        RECT 0.249 0.144 0.267 0.162 ;
        RECT 0.937 0.144 0.955 0.162 ;
        RECT 1.261 0.144 1.279 0.162 ;
        RECT 1.441 0.144 1.459 0.162 ;
        RECT 1.639 0.144 1.657 0.162 ;
        RECT 2.333 0.144 2.351 0.162 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.077 0.172 1.117 0.199 ;
        RECT 1.099 0.07 1.117 0.199 ;
        RECT 1.033 0.222 1.096 0.241 ;
        RECT 1.077 0.172 1.096 0.241 ;
      LAYER M2 ;
        RECT 0.983 0.216 1.238 0.234 ;
      LAYER V1 ;
        RECT 1.077 0.216 1.096 0.234 ;
    END
  END ENA
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.153 0.07 1.171 0.199 ;
      LAYER M2 ;
        RECT 0.983 0.072 1.238 0.09 ;
      LAYER V1 ;
        RECT 1.153 0.072 1.171 0.09 ;
    END
  END SE
  OBS
    LAYER M1 ;
      RECT 2.255 0.222 2.413 0.24 ;
      RECT 2.395 0.188 2.413 0.24 ;
      RECT 2.395 0.188 2.467 0.206 ;
      RECT 2.449 0.063 2.467 0.206 ;
      RECT 2.309 0.063 2.467 0.081 ;
      RECT 2.395 0.099 2.413 0.147 ;
      RECT 2.233 0.099 2.251 0.147 ;
      RECT 2.233 0.099 2.413 0.117 ;
      RECT 2.125 0.126 2.181 0.144 ;
      RECT 2.125 0.09 2.143 0.144 ;
      RECT 2.039 0.09 2.191 0.108 ;
      RECT 2.02 0.162 2.175 0.18 ;
      RECT 2.071 0.126 2.089 0.18 ;
      RECT 2.031 0.126 2.089 0.144 ;
      RECT 1.715 0.222 1.873 0.24 ;
      RECT 1.855 0.188 1.873 0.24 ;
      RECT 1.855 0.188 1.927 0.206 ;
      RECT 1.909 0.063 1.927 0.206 ;
      RECT 1.769 0.063 1.927 0.081 ;
      RECT 1.283 0.223 1.394 0.241 ;
      RECT 1.376 0.027 1.394 0.241 ;
      RECT 1.376 0.181 1.5 0.199 ;
      RECT 1.855 0.099 1.873 0.147 ;
      RECT 1.693 0.027 1.711 0.147 ;
      RECT 1.693 0.099 1.873 0.117 ;
      RECT 1.337 0.027 1.711 0.045 ;
      RECT 1.586 0.223 1.636 0.241 ;
      RECT 1.586 0.077 1.604 0.241 ;
      RECT 1.586 0.077 1.636 0.095 ;
      RECT 1.495 0.224 1.549 0.242 ;
      RECT 1.53 0.073 1.549 0.242 ;
      RECT 1.419 0.073 1.549 0.091 ;
      RECT 1.315 0.18 1.351 0.198 ;
      RECT 1.315 0.072 1.333 0.198 ;
      RECT 1.284 0.072 1.333 0.09 ;
      RECT 1.121 0.224 1.225 0.242 ;
      RECT 1.207 0.027 1.225 0.242 ;
      RECT 1.116 0.027 1.225 0.045 ;
      RECT 0.958 0.223 1.008 0.241 ;
      RECT 0.99 0.077 1.008 0.241 ;
      RECT 0.958 0.077 1.008 0.095 ;
      RECT 0.883 0.099 0.901 0.147 ;
      RECT 0.721 0.099 0.739 0.147 ;
      RECT 0.721 0.099 0.901 0.117 ;
      RECT 0.721 0.222 0.879 0.24 ;
      RECT 0.721 0.188 0.739 0.24 ;
      RECT 0.667 0.188 0.739 0.206 ;
      RECT 0.667 0.063 0.685 0.206 ;
      RECT 0.667 0.063 0.825 0.081 ;
      RECT 0.419 0.162 0.574 0.18 ;
      RECT 0.505 0.126 0.523 0.18 ;
      RECT 0.505 0.126 0.563 0.144 ;
      RECT 0.413 0.126 0.469 0.144 ;
      RECT 0.451 0.09 0.469 0.144 ;
      RECT 0.403 0.09 0.555 0.108 ;
      RECT 0.343 0.099 0.361 0.147 ;
      RECT 0.181 0.099 0.199 0.147 ;
      RECT 0.181 0.099 0.361 0.117 ;
      RECT 0.181 0.222 0.339 0.24 ;
      RECT 0.181 0.188 0.199 0.24 ;
      RECT 0.127 0.188 0.199 0.206 ;
      RECT 0.127 0.063 0.145 0.206 ;
      RECT 0.127 0.063 0.285 0.081 ;
    LAYER M2 ;
      RECT 0.337 0.108 2.257 0.126 ;
      RECT 0.983 0.18 1.609 0.198 ;
    LAYER V1 ;
      RECT 2.233 0.108 2.251 0.126 ;
      RECT 1.693 0.108 1.711 0.126 ;
      RECT 1.586 0.18 1.604 0.198 ;
      RECT 1.328 0.18 1.346 0.198 ;
      RECT 0.99 0.18 1.008 0.198 ;
      RECT 0.883 0.108 0.901 0.126 ;
      RECT 0.343 0.108 0.361 0.126 ;
  END
END ICGx4DC_ASAP7_75t_L

MACRO ICGx4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx4_ASAP7_75t_L 0 0 ;
  SIZE 1.134 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.199 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.89 0.225 1.062 0.243 ;
        RECT 1.044 0.027 1.062 0.243 ;
        RECT 0.889 0.027 1.062 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.199 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.134 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.134 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.229 0.144 0.635 0.162 ;
      LAYER M1 ;
        RECT 0.612 0.178 0.765 0.196 ;
        RECT 0.747 0.142 0.765 0.196 ;
        RECT 0.612 0.116 0.63 0.196 ;
        RECT 0.396 0.144 0.447 0.162 ;
        RECT 0.396 0.12 0.414 0.162 ;
        RECT 0.234 0.119 0.252 0.184 ;
      LAYER V1 ;
        RECT 0.234 0.144 0.252 0.162 ;
        RECT 0.414 0.144 0.432 0.162 ;
        RECT 0.612 0.144 0.63 0.162 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.688 0.222 0.846 0.24 ;
      RECT 0.828 0.188 0.846 0.24 ;
      RECT 0.828 0.188 0.9 0.206 ;
      RECT 0.882 0.063 0.9 0.206 ;
      RECT 0.742 0.063 0.9 0.081 ;
      RECT 0.256 0.223 0.367 0.241 ;
      RECT 0.349 0.027 0.367 0.241 ;
      RECT 0.349 0.181 0.473 0.199 ;
      RECT 0.828 0.099 0.846 0.147 ;
      RECT 0.666 0.027 0.684 0.147 ;
      RECT 0.666 0.099 0.846 0.117 ;
      RECT 0.31 0.027 0.684 0.045 ;
      RECT 0.559 0.223 0.609 0.241 ;
      RECT 0.559 0.077 0.577 0.241 ;
      RECT 0.559 0.077 0.609 0.095 ;
      RECT 0.468 0.224 0.522 0.242 ;
      RECT 0.503 0.073 0.522 0.242 ;
      RECT 0.392 0.073 0.522 0.091 ;
      RECT 0.288 0.18 0.324 0.198 ;
      RECT 0.288 0.072 0.306 0.198 ;
      RECT 0.257 0.072 0.306 0.09 ;
      RECT 0.037 0.224 0.198 0.242 ;
      RECT 0.18 0.027 0.198 0.242 ;
      RECT 0.089 0.027 0.198 0.045 ;
    LAYER M2 ;
      RECT 0.296 0.18 0.582 0.198 ;
    LAYER V1 ;
      RECT 0.559 0.18 0.577 0.198 ;
      RECT 0.301 0.18 0.319 0.198 ;
  END
END ICGx4_ASAP7_75t_L

MACRO ICGx5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx5_ASAP7_75t_L 0 0 ;
  SIZE 1.188 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.199 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.89 0.225 1.17 0.243 ;
        RECT 1.152 0.027 1.17 0.243 ;
        RECT 0.889 0.027 1.17 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.199 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.229 0.144 0.635 0.162 ;
      LAYER M1 ;
        RECT 0.612 0.178 0.765 0.196 ;
        RECT 0.747 0.142 0.765 0.196 ;
        RECT 0.612 0.116 0.63 0.196 ;
        RECT 0.396 0.144 0.447 0.162 ;
        RECT 0.396 0.12 0.414 0.162 ;
        RECT 0.234 0.119 0.252 0.184 ;
      LAYER V1 ;
        RECT 0.234 0.144 0.252 0.162 ;
        RECT 0.414 0.144 0.432 0.162 ;
        RECT 0.612 0.144 0.63 0.162 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.688 0.222 0.846 0.24 ;
      RECT 0.828 0.188 0.846 0.24 ;
      RECT 0.828 0.188 0.9 0.206 ;
      RECT 0.882 0.063 0.9 0.206 ;
      RECT 0.742 0.063 0.9 0.081 ;
      RECT 0.256 0.223 0.367 0.241 ;
      RECT 0.349 0.027 0.367 0.241 ;
      RECT 0.349 0.181 0.473 0.199 ;
      RECT 0.828 0.099 0.846 0.147 ;
      RECT 0.666 0.027 0.684 0.147 ;
      RECT 0.666 0.099 0.846 0.117 ;
      RECT 0.31 0.027 0.684 0.045 ;
      RECT 0.559 0.223 0.609 0.241 ;
      RECT 0.559 0.077 0.577 0.241 ;
      RECT 0.559 0.077 0.609 0.095 ;
      RECT 0.468 0.224 0.522 0.242 ;
      RECT 0.503 0.073 0.522 0.242 ;
      RECT 0.392 0.073 0.522 0.091 ;
      RECT 0.288 0.18 0.324 0.198 ;
      RECT 0.288 0.072 0.306 0.198 ;
      RECT 0.257 0.072 0.306 0.09 ;
      RECT 0.037 0.224 0.198 0.242 ;
      RECT 0.18 0.027 0.198 0.242 ;
      RECT 0.089 0.027 0.198 0.045 ;
    LAYER M2 ;
      RECT 0.296 0.18 0.582 0.198 ;
    LAYER V1 ;
      RECT 0.559 0.18 0.577 0.198 ;
      RECT 0.301 0.18 0.319 0.198 ;
  END
END ICGx5_ASAP7_75t_L

MACRO ICGx5p33DC_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx5p33DC_ASAP7_75t_L 0 0 ;
  SIZE 2.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.466 0.225 2.521 0.243 ;
        RECT 2.503 0.027 2.521 0.243 ;
        RECT 2.446 0.027 2.521 0.045 ;
        RECT 1.926 0.225 1.981 0.243 ;
        RECT 1.963 0.027 1.981 0.243 ;
        RECT 1.906 0.027 1.981 0.045 ;
        RECT 0.613 0.027 0.688 0.045 ;
        RECT 0.613 0.225 0.668 0.243 ;
        RECT 0.613 0.027 0.631 0.243 ;
        RECT 0.073 0.027 0.148 0.045 ;
        RECT 0.073 0.225 0.128 0.243 ;
        RECT 0.073 0.027 0.091 0.243 ;
      LAYER M2 ;
        RECT 0.062 0.036 2.532 0.054 ;
      LAYER V1 ;
        RECT 0.073 0.036 0.091 0.054 ;
        RECT 0.613 0.036 0.631 0.054 ;
        RECT 1.963 0.036 1.981 0.054 ;
        RECT 2.503 0.036 2.521 0.054 ;
    END
  END GCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.594 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 2.282 0.171 2.351 0.189 ;
        RECT 2.333 0.135 2.351 0.189 ;
        RECT 2.293 0.135 2.351 0.153 ;
        RECT 1.639 0.178 1.792 0.196 ;
        RECT 1.774 0.142 1.792 0.196 ;
        RECT 1.639 0.116 1.657 0.196 ;
        RECT 1.423 0.144 1.474 0.162 ;
        RECT 1.423 0.12 1.441 0.162 ;
        RECT 1.261 0.119 1.279 0.184 ;
        RECT 0.802 0.178 0.955 0.196 ;
        RECT 0.937 0.116 0.955 0.196 ;
        RECT 0.802 0.142 0.82 0.196 ;
        RECT 0.249 0.171 0.318 0.189 ;
        RECT 0.249 0.135 0.307 0.153 ;
        RECT 0.249 0.135 0.267 0.189 ;
      LAYER M2 ;
        RECT 0.236 0.144 2.359 0.162 ;
      LAYER V1 ;
        RECT 0.249 0.144 0.267 0.162 ;
        RECT 0.937 0.144 0.955 0.162 ;
        RECT 1.261 0.144 1.279 0.162 ;
        RECT 1.441 0.144 1.459 0.162 ;
        RECT 1.639 0.144 1.657 0.162 ;
        RECT 2.333 0.144 2.351 0.162 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.077 0.172 1.117 0.199 ;
        RECT 1.099 0.07 1.117 0.199 ;
        RECT 1.033 0.222 1.096 0.241 ;
        RECT 1.077 0.172 1.096 0.241 ;
      LAYER M2 ;
        RECT 0.983 0.216 1.238 0.234 ;
      LAYER V1 ;
        RECT 1.077 0.216 1.096 0.234 ;
    END
  END ENA
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.153 0.07 1.171 0.199 ;
      LAYER M2 ;
        RECT 0.983 0.072 1.238 0.09 ;
      LAYER V1 ;
        RECT 1.153 0.072 1.171 0.09 ;
    END
  END SE
  OBS
    LAYER M1 ;
      RECT 2.255 0.222 2.413 0.24 ;
      RECT 2.395 0.188 2.413 0.24 ;
      RECT 2.395 0.188 2.467 0.206 ;
      RECT 2.449 0.063 2.467 0.206 ;
      RECT 2.309 0.063 2.467 0.081 ;
      RECT 2.395 0.099 2.413 0.147 ;
      RECT 2.233 0.099 2.251 0.147 ;
      RECT 2.233 0.099 2.413 0.117 ;
      RECT 2.125 0.126 2.181 0.144 ;
      RECT 2.125 0.09 2.143 0.144 ;
      RECT 2.039 0.09 2.191 0.108 ;
      RECT 2.02 0.162 2.175 0.18 ;
      RECT 2.071 0.126 2.089 0.18 ;
      RECT 2.031 0.126 2.089 0.144 ;
      RECT 1.715 0.222 1.873 0.24 ;
      RECT 1.855 0.188 1.873 0.24 ;
      RECT 1.855 0.188 1.927 0.206 ;
      RECT 1.909 0.063 1.927 0.206 ;
      RECT 1.769 0.063 1.927 0.081 ;
      RECT 1.283 0.223 1.394 0.241 ;
      RECT 1.376 0.027 1.394 0.241 ;
      RECT 1.376 0.181 1.5 0.199 ;
      RECT 1.855 0.099 1.873 0.147 ;
      RECT 1.693 0.027 1.711 0.147 ;
      RECT 1.693 0.099 1.873 0.117 ;
      RECT 1.337 0.027 1.711 0.045 ;
      RECT 1.586 0.223 1.636 0.241 ;
      RECT 1.586 0.077 1.604 0.241 ;
      RECT 1.586 0.077 1.636 0.095 ;
      RECT 1.495 0.224 1.549 0.242 ;
      RECT 1.53 0.073 1.549 0.242 ;
      RECT 1.419 0.073 1.549 0.091 ;
      RECT 1.315 0.18 1.351 0.198 ;
      RECT 1.315 0.072 1.333 0.198 ;
      RECT 1.284 0.072 1.333 0.09 ;
      RECT 1.121 0.224 1.225 0.242 ;
      RECT 1.207 0.027 1.225 0.242 ;
      RECT 1.116 0.027 1.225 0.045 ;
      RECT 0.958 0.223 1.008 0.241 ;
      RECT 0.99 0.077 1.008 0.241 ;
      RECT 0.958 0.077 1.008 0.095 ;
      RECT 0.883 0.099 0.901 0.147 ;
      RECT 0.721 0.099 0.739 0.147 ;
      RECT 0.721 0.099 0.901 0.117 ;
      RECT 0.721 0.222 0.879 0.24 ;
      RECT 0.721 0.188 0.739 0.24 ;
      RECT 0.667 0.188 0.739 0.206 ;
      RECT 0.667 0.063 0.685 0.206 ;
      RECT 0.667 0.063 0.825 0.081 ;
      RECT 0.419 0.162 0.574 0.18 ;
      RECT 0.505 0.126 0.523 0.18 ;
      RECT 0.505 0.126 0.563 0.144 ;
      RECT 0.413 0.126 0.469 0.144 ;
      RECT 0.451 0.09 0.469 0.144 ;
      RECT 0.403 0.09 0.555 0.108 ;
      RECT 0.343 0.099 0.361 0.147 ;
      RECT 0.181 0.099 0.199 0.147 ;
      RECT 0.181 0.099 0.361 0.117 ;
      RECT 0.181 0.222 0.339 0.24 ;
      RECT 0.181 0.188 0.199 0.24 ;
      RECT 0.127 0.188 0.199 0.206 ;
      RECT 0.127 0.063 0.145 0.206 ;
      RECT 0.127 0.063 0.285 0.081 ;
    LAYER M2 ;
      RECT 0.337 0.108 2.257 0.126 ;
      RECT 0.983 0.18 1.609 0.198 ;
    LAYER V1 ;
      RECT 2.233 0.108 2.251 0.126 ;
      RECT 1.693 0.108 1.711 0.126 ;
      RECT 1.586 0.18 1.604 0.198 ;
      RECT 1.328 0.18 1.346 0.198 ;
      RECT 0.99 0.18 1.008 0.198 ;
      RECT 0.883 0.108 0.901 0.126 ;
      RECT 0.343 0.108 0.361 0.126 ;
  END
END ICGx5p33DC_ASAP7_75t_L

MACRO ICGx6p67DC_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx6p67DC_ASAP7_75t_L 0 0 ;
  SIZE 2.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.466 0.225 2.521 0.243 ;
        RECT 2.503 0.027 2.521 0.243 ;
        RECT 2.446 0.027 2.521 0.045 ;
        RECT 1.926 0.225 1.981 0.243 ;
        RECT 1.963 0.027 1.981 0.243 ;
        RECT 1.906 0.027 1.981 0.045 ;
        RECT 0.613 0.027 0.688 0.045 ;
        RECT 0.613 0.225 0.668 0.243 ;
        RECT 0.613 0.027 0.631 0.243 ;
        RECT 0.073 0.027 0.148 0.045 ;
        RECT 0.073 0.225 0.128 0.243 ;
        RECT 0.073 0.027 0.091 0.243 ;
      LAYER M2 ;
        RECT 0.062 0.036 2.532 0.054 ;
      LAYER V1 ;
        RECT 0.073 0.036 0.091 0.054 ;
        RECT 0.613 0.036 0.631 0.054 ;
        RECT 1.963 0.036 1.981 0.054 ;
        RECT 2.503 0.036 2.521 0.054 ;
    END
  END GCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.594 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 2.282 0.171 2.351 0.189 ;
        RECT 2.333 0.135 2.351 0.189 ;
        RECT 2.293 0.135 2.351 0.153 ;
        RECT 1.639 0.178 1.792 0.196 ;
        RECT 1.774 0.142 1.792 0.196 ;
        RECT 1.639 0.116 1.657 0.196 ;
        RECT 1.423 0.144 1.474 0.162 ;
        RECT 1.423 0.12 1.441 0.162 ;
        RECT 1.261 0.119 1.279 0.184 ;
        RECT 0.802 0.178 0.955 0.196 ;
        RECT 0.937 0.116 0.955 0.196 ;
        RECT 0.802 0.142 0.82 0.196 ;
        RECT 0.249 0.171 0.318 0.189 ;
        RECT 0.249 0.135 0.307 0.153 ;
        RECT 0.249 0.135 0.267 0.189 ;
      LAYER M2 ;
        RECT 0.236 0.144 2.359 0.162 ;
      LAYER V1 ;
        RECT 0.249 0.144 0.267 0.162 ;
        RECT 0.937 0.144 0.955 0.162 ;
        RECT 1.261 0.144 1.279 0.162 ;
        RECT 1.441 0.144 1.459 0.162 ;
        RECT 1.639 0.144 1.657 0.162 ;
        RECT 2.333 0.144 2.351 0.162 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.077 0.172 1.117 0.199 ;
        RECT 1.099 0.07 1.117 0.199 ;
        RECT 1.033 0.222 1.096 0.241 ;
        RECT 1.077 0.172 1.096 0.241 ;
      LAYER M2 ;
        RECT 0.983 0.216 1.238 0.234 ;
      LAYER V1 ;
        RECT 1.077 0.216 1.096 0.234 ;
    END
  END ENA
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.153 0.07 1.171 0.199 ;
      LAYER M2 ;
        RECT 0.983 0.072 1.238 0.09 ;
      LAYER V1 ;
        RECT 1.153 0.072 1.171 0.09 ;
    END
  END SE
  OBS
    LAYER M1 ;
      RECT 2.255 0.222 2.413 0.24 ;
      RECT 2.395 0.188 2.413 0.24 ;
      RECT 2.395 0.188 2.467 0.206 ;
      RECT 2.449 0.063 2.467 0.206 ;
      RECT 2.309 0.063 2.467 0.081 ;
      RECT 2.395 0.099 2.413 0.147 ;
      RECT 2.233 0.099 2.251 0.147 ;
      RECT 2.233 0.099 2.413 0.117 ;
      RECT 2.125 0.126 2.181 0.144 ;
      RECT 2.125 0.09 2.143 0.144 ;
      RECT 2.039 0.09 2.191 0.108 ;
      RECT 2.02 0.162 2.175 0.18 ;
      RECT 2.071 0.126 2.089 0.18 ;
      RECT 2.031 0.126 2.089 0.144 ;
      RECT 1.715 0.222 1.873 0.24 ;
      RECT 1.855 0.188 1.873 0.24 ;
      RECT 1.855 0.188 1.927 0.206 ;
      RECT 1.909 0.063 1.927 0.206 ;
      RECT 1.769 0.063 1.927 0.081 ;
      RECT 1.283 0.223 1.394 0.241 ;
      RECT 1.376 0.027 1.394 0.241 ;
      RECT 1.376 0.181 1.5 0.199 ;
      RECT 1.855 0.099 1.873 0.147 ;
      RECT 1.693 0.027 1.711 0.147 ;
      RECT 1.693 0.099 1.873 0.117 ;
      RECT 1.337 0.027 1.711 0.045 ;
      RECT 1.586 0.223 1.636 0.241 ;
      RECT 1.586 0.077 1.604 0.241 ;
      RECT 1.586 0.077 1.636 0.095 ;
      RECT 1.495 0.224 1.549 0.242 ;
      RECT 1.53 0.073 1.549 0.242 ;
      RECT 1.419 0.073 1.549 0.091 ;
      RECT 1.315 0.18 1.351 0.198 ;
      RECT 1.315 0.072 1.333 0.198 ;
      RECT 1.284 0.072 1.333 0.09 ;
      RECT 1.121 0.224 1.225 0.242 ;
      RECT 1.207 0.027 1.225 0.242 ;
      RECT 1.116 0.027 1.225 0.045 ;
      RECT 0.958 0.223 1.008 0.241 ;
      RECT 0.99 0.077 1.008 0.241 ;
      RECT 0.958 0.077 1.008 0.095 ;
      RECT 0.883 0.099 0.901 0.147 ;
      RECT 0.721 0.099 0.739 0.147 ;
      RECT 0.721 0.099 0.901 0.117 ;
      RECT 0.721 0.222 0.879 0.24 ;
      RECT 0.721 0.188 0.739 0.24 ;
      RECT 0.667 0.188 0.739 0.206 ;
      RECT 0.667 0.063 0.685 0.206 ;
      RECT 0.667 0.063 0.825 0.081 ;
      RECT 0.419 0.162 0.574 0.18 ;
      RECT 0.505 0.126 0.523 0.18 ;
      RECT 0.505 0.126 0.563 0.144 ;
      RECT 0.413 0.126 0.469 0.144 ;
      RECT 0.451 0.09 0.469 0.144 ;
      RECT 0.403 0.09 0.555 0.108 ;
      RECT 0.343 0.099 0.361 0.147 ;
      RECT 0.181 0.099 0.199 0.147 ;
      RECT 0.181 0.099 0.361 0.117 ;
      RECT 0.181 0.222 0.339 0.24 ;
      RECT 0.181 0.188 0.199 0.24 ;
      RECT 0.127 0.188 0.199 0.206 ;
      RECT 0.127 0.063 0.145 0.206 ;
      RECT 0.127 0.063 0.285 0.081 ;
    LAYER M2 ;
      RECT 0.337 0.108 2.257 0.126 ;
      RECT 0.983 0.18 1.609 0.198 ;
    LAYER V1 ;
      RECT 2.233 0.108 2.251 0.126 ;
      RECT 1.693 0.108 1.711 0.126 ;
      RECT 1.586 0.18 1.604 0.198 ;
      RECT 1.328 0.18 1.346 0.198 ;
      RECT 0.99 0.18 1.008 0.198 ;
      RECT 0.883 0.108 0.901 0.126 ;
      RECT 0.343 0.108 0.361 0.126 ;
  END
END ICGx6p67DC_ASAP7_75t_L

MACRO ICGx8DC_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx8DC_ASAP7_75t_L 0 0 ;
  SIZE 2.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.466 0.225 2.521 0.243 ;
        RECT 2.503 0.027 2.521 0.243 ;
        RECT 2.446 0.027 2.521 0.045 ;
        RECT 1.926 0.225 1.981 0.243 ;
        RECT 1.963 0.027 1.981 0.243 ;
        RECT 1.906 0.027 1.981 0.045 ;
        RECT 0.613 0.027 0.688 0.045 ;
        RECT 0.613 0.225 0.668 0.243 ;
        RECT 0.613 0.027 0.631 0.243 ;
        RECT 0.073 0.027 0.148 0.045 ;
        RECT 0.073 0.225 0.128 0.243 ;
        RECT 0.073 0.027 0.091 0.243 ;
      LAYER M2 ;
        RECT 0.062 0.036 2.532 0.054 ;
      LAYER V1 ;
        RECT 0.073 0.036 0.091 0.054 ;
        RECT 0.613 0.036 0.631 0.054 ;
        RECT 1.963 0.036 1.981 0.054 ;
        RECT 2.503 0.036 2.521 0.054 ;
    END
  END GCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.594 0.009 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 2.282 0.171 2.351 0.189 ;
        RECT 2.333 0.135 2.351 0.189 ;
        RECT 2.293 0.135 2.351 0.153 ;
        RECT 1.639 0.178 1.792 0.196 ;
        RECT 1.774 0.142 1.792 0.196 ;
        RECT 1.639 0.116 1.657 0.196 ;
        RECT 1.423 0.144 1.474 0.162 ;
        RECT 1.423 0.12 1.441 0.162 ;
        RECT 1.261 0.119 1.279 0.184 ;
        RECT 0.802 0.178 0.955 0.196 ;
        RECT 0.937 0.116 0.955 0.196 ;
        RECT 0.802 0.142 0.82 0.196 ;
        RECT 0.249 0.171 0.318 0.189 ;
        RECT 0.249 0.135 0.307 0.153 ;
        RECT 0.249 0.135 0.267 0.189 ;
      LAYER M2 ;
        RECT 0.236 0.144 2.359 0.162 ;
      LAYER V1 ;
        RECT 0.249 0.144 0.267 0.162 ;
        RECT 0.937 0.144 0.955 0.162 ;
        RECT 1.261 0.144 1.279 0.162 ;
        RECT 1.441 0.144 1.459 0.162 ;
        RECT 1.639 0.144 1.657 0.162 ;
        RECT 2.333 0.144 2.351 0.162 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.077 0.172 1.117 0.199 ;
        RECT 1.099 0.07 1.117 0.199 ;
        RECT 1.033 0.222 1.096 0.241 ;
        RECT 1.077 0.172 1.096 0.241 ;
      LAYER M2 ;
        RECT 0.983 0.216 1.238 0.234 ;
      LAYER V1 ;
        RECT 1.077 0.216 1.096 0.234 ;
    END
  END ENA
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.153 0.07 1.171 0.199 ;
      LAYER M2 ;
        RECT 0.983 0.072 1.238 0.09 ;
      LAYER V1 ;
        RECT 1.153 0.072 1.171 0.09 ;
    END
  END SE
  OBS
    LAYER M1 ;
      RECT 2.255 0.222 2.413 0.24 ;
      RECT 2.395 0.188 2.413 0.24 ;
      RECT 2.395 0.188 2.467 0.206 ;
      RECT 2.449 0.063 2.467 0.206 ;
      RECT 2.309 0.063 2.467 0.081 ;
      RECT 2.395 0.099 2.413 0.147 ;
      RECT 2.233 0.099 2.251 0.147 ;
      RECT 2.233 0.099 2.413 0.117 ;
      RECT 2.125 0.126 2.181 0.144 ;
      RECT 2.125 0.09 2.143 0.144 ;
      RECT 2.039 0.09 2.191 0.108 ;
      RECT 2.02 0.162 2.175 0.18 ;
      RECT 2.071 0.126 2.089 0.18 ;
      RECT 2.031 0.126 2.089 0.144 ;
      RECT 1.715 0.222 1.873 0.24 ;
      RECT 1.855 0.188 1.873 0.24 ;
      RECT 1.855 0.188 1.927 0.206 ;
      RECT 1.909 0.063 1.927 0.206 ;
      RECT 1.769 0.063 1.927 0.081 ;
      RECT 1.283 0.223 1.394 0.241 ;
      RECT 1.376 0.027 1.394 0.241 ;
      RECT 1.376 0.181 1.5 0.199 ;
      RECT 1.855 0.099 1.873 0.147 ;
      RECT 1.693 0.027 1.711 0.147 ;
      RECT 1.693 0.099 1.873 0.117 ;
      RECT 1.337 0.027 1.711 0.045 ;
      RECT 1.586 0.223 1.636 0.241 ;
      RECT 1.586 0.077 1.604 0.241 ;
      RECT 1.586 0.077 1.636 0.095 ;
      RECT 1.495 0.224 1.549 0.242 ;
      RECT 1.53 0.073 1.549 0.242 ;
      RECT 1.419 0.073 1.549 0.091 ;
      RECT 1.315 0.18 1.351 0.198 ;
      RECT 1.315 0.072 1.333 0.198 ;
      RECT 1.284 0.072 1.333 0.09 ;
      RECT 1.121 0.224 1.225 0.242 ;
      RECT 1.207 0.027 1.225 0.242 ;
      RECT 1.116 0.027 1.225 0.045 ;
      RECT 0.958 0.223 1.008 0.241 ;
      RECT 0.99 0.077 1.008 0.241 ;
      RECT 0.958 0.077 1.008 0.095 ;
      RECT 0.883 0.099 0.901 0.147 ;
      RECT 0.721 0.099 0.739 0.147 ;
      RECT 0.721 0.099 0.901 0.117 ;
      RECT 0.721 0.222 0.879 0.24 ;
      RECT 0.721 0.188 0.739 0.24 ;
      RECT 0.667 0.188 0.739 0.206 ;
      RECT 0.667 0.063 0.685 0.206 ;
      RECT 0.667 0.063 0.825 0.081 ;
      RECT 0.419 0.162 0.574 0.18 ;
      RECT 0.505 0.126 0.523 0.18 ;
      RECT 0.505 0.126 0.563 0.144 ;
      RECT 0.413 0.126 0.469 0.144 ;
      RECT 0.451 0.09 0.469 0.144 ;
      RECT 0.403 0.09 0.555 0.108 ;
      RECT 0.343 0.099 0.361 0.147 ;
      RECT 0.181 0.099 0.199 0.147 ;
      RECT 0.181 0.099 0.361 0.117 ;
      RECT 0.181 0.222 0.339 0.24 ;
      RECT 0.181 0.188 0.199 0.24 ;
      RECT 0.127 0.188 0.199 0.206 ;
      RECT 0.127 0.063 0.145 0.206 ;
      RECT 0.127 0.063 0.285 0.081 ;
    LAYER M2 ;
      RECT 0.337 0.108 2.257 0.126 ;
      RECT 0.983 0.18 1.609 0.198 ;
    LAYER V1 ;
      RECT 2.233 0.108 2.251 0.126 ;
      RECT 1.693 0.108 1.711 0.126 ;
      RECT 1.586 0.18 1.604 0.198 ;
      RECT 1.328 0.18 1.346 0.198 ;
      RECT 0.99 0.18 1.008 0.198 ;
      RECT 0.883 0.108 0.901 0.126 ;
      RECT 0.343 0.108 0.361 0.126 ;
  END
END ICGx8DC_ASAP7_75t_L

MACRO INVx11_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx11_ASAP7_75t_L 0 0 ;
  SIZE 0.702 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.702 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.684 0.243 ;
        RECT 0.666 0.027 0.684 0.243 ;
        RECT 0.094 0.027 0.684 0.045 ;
    END
  END Y
END INVx11_ASAP7_75t_L

MACRO INVx13_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx13_ASAP7_75t_L 0 0 ;
  SIZE 0.81 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.81 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.792 0.243 ;
        RECT 0.774 0.027 0.792 0.243 ;
        RECT 0.094 0.027 0.792 0.045 ;
    END
  END Y
END INVx13_ASAP7_75t_L

MACRO INVx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx1_ASAP7_75t_L 0 0 ;
  SIZE 0.162 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.162 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.144 0.243 ;
        RECT 0.126 0.027 0.144 0.243 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END Y
END INVx1_ASAP7_75t_L

MACRO INVx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx2_ASAP7_75t_L 0 0 ;
  SIZE 0.216 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.216 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.144 0.243 ;
        RECT 0.126 0.027 0.144 0.243 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END Y
END INVx2_ASAP7_75t_L

MACRO INVx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx3_ASAP7_75t_L 0 0 ;
  SIZE 0.27 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.27 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.252 0.243 ;
        RECT 0.234 0.027 0.252 0.243 ;
        RECT 0.094 0.027 0.252 0.045 ;
    END
  END Y
END INVx3_ASAP7_75t_L

MACRO INVx4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx4_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.306 0.243 ;
        RECT 0.288 0.027 0.306 0.243 ;
        RECT 0.094 0.027 0.306 0.045 ;
    END
  END Y
END INVx4_ASAP7_75t_L

MACRO INVx5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx5_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.36 0.243 ;
        RECT 0.342 0.027 0.36 0.243 ;
        RECT 0.094 0.027 0.36 0.045 ;
    END
  END Y
END INVx5_ASAP7_75t_L

MACRO INVx6_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx6_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.094 0.027 0.414 0.045 ;
    END
  END Y
END INVx6_ASAP7_75t_L

MACRO INVx8_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx8_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.522 0.243 ;
        RECT 0.504 0.027 0.522 0.243 ;
        RECT 0.094 0.027 0.522 0.045 ;
    END
  END Y
END INVx8_ASAP7_75t_L

MACRO INVxp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVxp33_ASAP7_75t_L 0 0 ;
  SIZE 0.162 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.162 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.144 0.243 ;
        RECT 0.126 0.027 0.144 0.243 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END Y
END INVxp33_ASAP7_75t_L

MACRO INVxp67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVxp67_ASAP7_75t_L 0 0 ;
  SIZE 0.162 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.162 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.144 0.243 ;
        RECT 0.126 0.027 0.144 0.243 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END Y
END INVxp67_ASAP7_75t_L

MACRO MAJIxp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJIxp5_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.164 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.126 0.257 0.144 ;
        RECT 0.018 0.189 0.198 0.207 ;
        RECT 0.18 0.126 0.198 0.207 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.034 0.036 0.207 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.255 0.189 0.361 0.207 ;
        RECT 0.343 0.063 0.361 0.207 ;
        RECT 0.255 0.063 0.361 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.027 0.338 0.045 ;
      RECT 0.094 0.225 0.338 0.243 ;
  END
END MAJIxp5_ASAP7_75t_L

MACRO MAJx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJx2_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.164 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.189 0.333 0.207 ;
        RECT 0.315 0.106 0.333 0.207 ;
        RECT 0.283 0.126 0.333 0.144 ;
        RECT 0.18 0.126 0.198 0.207 ;
        RECT 0.121 0.126 0.198 0.144 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.364 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.189 0.123 0.207 ;
      RECT 0.018 0.063 0.036 0.207 ;
      RECT 0.368 0.063 0.386 0.149 ;
      RECT 0.018 0.063 0.386 0.081 ;
      RECT 0.04 0.027 0.284 0.045 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END MAJx2_ASAP7_75t_L

MACRO MAJx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJx3_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.164 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.189 0.333 0.207 ;
        RECT 0.315 0.106 0.333 0.207 ;
        RECT 0.283 0.126 0.333 0.144 ;
        RECT 0.18 0.126 0.198 0.207 ;
        RECT 0.121 0.126 0.198 0.144 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.225 0.504 0.243 ;
        RECT 0.364 0.027 0.504 0.045 ;
        RECT 0.45 0.027 0.468 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.189 0.123 0.207 ;
      RECT 0.018 0.063 0.036 0.207 ;
      RECT 0.368 0.063 0.386 0.149 ;
      RECT 0.018 0.063 0.386 0.081 ;
      RECT 0.04 0.027 0.284 0.045 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END MAJx3_ASAP7_75t_L

MACRO NAND2x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.084 0.144 ;
        RECT 0.018 0.065 0.036 0.236 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.306 0.243 ;
        RECT 0.288 0.063 0.306 0.243 ;
        RECT 0.202 0.063 0.306 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.284 0.045 ;
  END
END NAND2x1_ASAP7_75t_L

MACRO NAND2x1p5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1p5_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.084 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.126 0.257 0.144 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.261 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.063 0.338 0.081 ;
      RECT 0.094 0.027 0.225 0.045 ;
  END
END NAND2x1p5_ASAP7_75t_L

MACRO NAND2x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x2_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.189 0.279 0.207 ;
        RECT 0.261 0.106 0.279 0.207 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.099 0.468 0.177 ;
        RECT 0.322 0.099 0.468 0.117 ;
        RECT 0.322 0.063 0.34 0.117 ;
        RECT 0.2 0.063 0.34 0.081 ;
        RECT 0.072 0.099 0.218 0.117 ;
        RECT 0.2 0.063 0.218 0.117 ;
        RECT 0.072 0.189 0.109 0.207 ;
        RECT 0.072 0.099 0.09 0.207 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.522 0.243 ;
        RECT 0.504 0.063 0.522 0.243 ;
        RECT 0.418 0.063 0.522 0.081 ;
        RECT 0.018 0.063 0.122 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.5 0.045 ;
  END
END NAND2x2_ASAP7_75t_L

MACRO NAND2xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.216 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.216 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.198 0.243 ;
        RECT 0.18 0.027 0.198 0.243 ;
        RECT 0.143 0.027 0.198 0.045 ;
    END
  END Y
END NAND2xp33_ASAP7_75t_L

MACRO NAND2xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.216 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.106 0.063 0.144 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.216 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.198 0.243 ;
        RECT 0.18 0.027 0.198 0.243 ;
        RECT 0.143 0.027 0.198 0.045 ;
    END
  END Y
END NAND2xp5_ASAP7_75t_L

MACRO NAND2xp67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp67_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.125 0.095 0.143 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.215 0.189 0.252 0.207 ;
        RECT 0.234 0.106 0.252 0.207 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.225 0.306 0.243 ;
        RECT 0.288 0.063 0.306 0.243 ;
        RECT 0.202 0.063 0.306 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.284 0.045 ;
  END
END NAND2xp67_ASAP7_75t_L

MACRO NAND3x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x1_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.402 0.18 0.468 0.198 ;
        RECT 0.45 0.108 0.468 0.198 ;
        RECT 0.4 0.108 0.468 0.126 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.243 0.18 0.306 0.198 ;
        RECT 0.288 0.108 0.306 0.198 ;
        RECT 0.246 0.108 0.306 0.126 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.061 0.103 0.079 0.203 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.225 0.576 0.243 ;
        RECT 0.558 0.063 0.576 0.243 ;
        RECT 0.418 0.063 0.576 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.256 0.027 0.5 0.045 ;
      RECT 0.094 0.063 0.338 0.081 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END NAND3x1_ASAP7_75t_L

MACRO NAND3x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x2_ASAP7_75t_L 0 0 ;
  SIZE 1.08 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.189 0.743 0.207 ;
        RECT 0.725 0.106 0.743 0.207 ;
        RECT 0.338 0.106 0.356 0.207 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.547 0.106 0.565 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.08 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 1.062 0.243 ;
        RECT 1.044 0.063 1.062 0.243 ;
        RECT 0.904 0.063 1.062 0.081 ;
        RECT 0.018 0.063 0.176 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.169 0.18 0.908 0.198 ;
      LAYER M1 ;
        RECT 0.866 0.189 0.903 0.207 ;
        RECT 0.885 0.108 0.903 0.207 ;
        RECT 0.174 0.189 0.211 0.207 ;
        RECT 0.174 0.106 0.192 0.207 ;
      LAYER V1 ;
        RECT 0.174 0.18 0.192 0.198 ;
        RECT 0.885 0.18 0.903 0.198 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 0.742 0.027 0.986 0.045 ;
      RECT 0.256 0.063 0.824 0.081 ;
      RECT 0.418 0.027 0.662 0.045 ;
      RECT 0.094 0.027 0.338 0.045 ;
  END
END NAND3x2_ASAP7_75t_L

MACRO NAND3xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.27 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.034 0.198 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.27 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.176 0.243 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
END NAND3xp33_ASAP7_75t_L

MACRO NAND4xp25_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4xp25_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.034 0.198 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.2 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.034 0.09 0.2 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.04 0.225 0.306 0.243 ;
        RECT 0.288 0.027 0.306 0.243 ;
        RECT 0.256 0.027 0.306 0.045 ;
    END
  END Y
END NAND4xp25_ASAP7_75t_L

MACRO NAND4xp75_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4xp75_ASAP7_75t_L 0 0 ;
  SIZE 0.756 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.106 0.63 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.101 0.549 0.119 ;
        RECT 0.531 0.07 0.549 0.119 ;
        RECT 0.504 0.101 0.522 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.101 0.306 0.2 ;
        RECT 0.207 0.101 0.306 0.119 ;
        RECT 0.207 0.07 0.225 0.119 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.225 0.057 0.243 ;
        RECT 0.018 0.027 0.057 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.756 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.738 0.243 ;
        RECT 0.72 0.063 0.738 0.243 ;
        RECT 0.58 0.063 0.738 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.412 0.027 0.666 0.045 ;
      RECT 0.256 0.063 0.499 0.081 ;
      RECT 0.092 0.027 0.34 0.045 ;
  END
END NAND4xp75_ASAP7_75t_L

MACRO NAND5xp2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND5xp2_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.034 0.144 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.034 0.198 0.2 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.034 0.252 0.2 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.034 0.306 0.2 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.009 0.225 0.317 0.243 ;
        RECT 0.009 0.027 0.07 0.045 ;
        RECT 0.009 0.027 0.027 0.243 ;
    END
  END Y
END NAND5xp2_ASAP7_75t_L

MACRO NOR2x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.084 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.126 0.23 0.144 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.189 0.306 0.207 ;
        RECT 0.288 0.027 0.306 0.207 ;
        RECT 0.094 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END NOR2x1_ASAP7_75t_L

MACRO NOR2x1p5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1p5_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.084 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.126 0.257 0.144 ;
        RECT 0.126 0.063 0.163 0.081 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.094 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.189 0.338 0.207 ;
      RECT 0.094 0.225 0.225 0.243 ;
  END
END NOR2x1p5_ASAP7_75t_L

MACRO NOR2x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x2_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.063 0.279 0.164 ;
        RECT 0.242 0.063 0.279 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.322 0.153 0.468 0.171 ;
        RECT 0.45 0.093 0.468 0.171 ;
        RECT 0.2 0.189 0.34 0.207 ;
        RECT 0.322 0.153 0.34 0.207 ;
        RECT 0.2 0.153 0.218 0.207 ;
        RECT 0.072 0.153 0.218 0.171 ;
        RECT 0.072 0.063 0.109 0.081 ;
        RECT 0.072 0.063 0.09 0.171 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.189 0.522 0.207 ;
        RECT 0.504 0.027 0.522 0.207 ;
        RECT 0.018 0.027 0.522 0.045 ;
        RECT 0.018 0.189 0.122 0.207 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.5 0.243 ;
  END
END NOR2x2_ASAP7_75t_L

MACRO NOR2xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.216 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.225 0.055 0.243 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.216 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.143 0.225 0.198 0.243 ;
        RECT 0.18 0.027 0.198 0.243 ;
        RECT 0.094 0.027 0.198 0.045 ;
    END
  END Y
END NOR2xp33_ASAP7_75t_L

MACRO NOR2xp67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2xp67_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.127 0.095 0.145 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.126 0.257 0.144 ;
        RECT 0.126 0.063 0.163 0.081 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.189 0.306 0.207 ;
        RECT 0.288 0.027 0.306 0.207 ;
        RECT 0.148 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END NOR2xp67_ASAP7_75t_L

MACRO NOR3x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x1_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.153 0.468 0.171 ;
        RECT 0.45 0.063 0.468 0.171 ;
        RECT 0.396 0.063 0.468 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.153 0.306 0.171 ;
        RECT 0.288 0.063 0.306 0.171 ;
        RECT 0.234 0.063 0.306 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.09 0.144 ;
        RECT 0.018 0.189 0.055 0.207 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.189 0.576 0.207 ;
        RECT 0.558 0.027 0.576 0.207 ;
        RECT 0.202 0.027 0.576 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.256 0.225 0.5 0.243 ;
      RECT 0.094 0.189 0.338 0.207 ;
      RECT 0.04 0.225 0.176 0.243 ;
  END
END NOR3x1_ASAP7_75t_L

MACRO NOR3x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x2_ASAP7_75t_L 0 0 ;
  SIZE 1.08 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.725 0.063 0.743 0.164 ;
        RECT 0.338 0.063 0.743 0.081 ;
        RECT 0.338 0.063 0.356 0.164 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.547 0.106 0.565 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.08 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.904 0.189 1.062 0.207 ;
        RECT 1.044 0.027 1.062 0.207 ;
        RECT 0.018 0.027 1.062 0.045 ;
        RECT 0.018 0.189 0.176 0.207 ;
        RECT 0.018 0.027 0.036 0.207 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.169 0.072 0.908 0.09 ;
      LAYER M1 ;
        RECT 0.885 0.063 0.903 0.162 ;
        RECT 0.866 0.063 0.903 0.081 ;
        RECT 0.174 0.063 0.211 0.081 ;
        RECT 0.174 0.063 0.192 0.164 ;
      LAYER V1 ;
        RECT 0.174 0.072 0.192 0.09 ;
        RECT 0.885 0.072 0.903 0.09 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 0.742 0.225 0.986 0.243 ;
      RECT 0.256 0.189 0.824 0.207 ;
      RECT 0.418 0.225 0.662 0.243 ;
      RECT 0.094 0.225 0.338 0.243 ;
  END
END NOR3x2_ASAP7_75t_L

MACRO NOR3xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.27 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.236 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.236 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.27 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.176 0.045 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
END NOR3xp33_ASAP7_75t_L

MACRO NOR4xp25_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4xp25_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.236 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.236 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.236 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.225 0.306 0.243 ;
        RECT 0.288 0.027 0.306 0.243 ;
        RECT 0.04 0.027 0.306 0.045 ;
    END
  END Y
END NOR4xp25_ASAP7_75t_L

MACRO NOR4xp75_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4xp75_ASAP7_75t_L 0 0 ;
  SIZE 0.756 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.07 0.63 0.164 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.531 0.151 0.549 0.2 ;
        RECT 0.504 0.151 0.549 0.169 ;
        RECT 0.504 0.07 0.522 0.169 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.151 0.306 0.169 ;
        RECT 0.288 0.07 0.306 0.169 ;
        RECT 0.207 0.151 0.225 0.2 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.225 0.057 0.243 ;
        RECT 0.018 0.027 0.057 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.756 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.189 0.738 0.207 ;
        RECT 0.72 0.027 0.738 0.207 ;
        RECT 0.094 0.027 0.738 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.412 0.225 0.666 0.243 ;
      RECT 0.256 0.189 0.499 0.207 ;
      RECT 0.092 0.225 0.34 0.243 ;
  END
END NOR4xp75_ASAP7_75t_L

MACRO NOR5xp2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR5xp2_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.198 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.236 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.236 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.236 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.236 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.027 0.338 0.045 ;
        RECT 0.017 0.225 0.07 0.243 ;
        RECT 0.017 0.027 0.037 0.243 ;
    END
  END Y
END NOR5xp2_ASAP7_75t_L

MACRO O2A1O1Ixp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN O2A1O1Ixp33_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.2 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.206 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.225 0.306 0.243 ;
        RECT 0.288 0.027 0.306 0.243 ;
        RECT 0.094 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.225 0.243 ;
      RECT 0.04 0.063 0.176 0.081 ;
  END
END O2A1O1Ixp33_ASAP7_75t_L

MACRO O2A1O1Ixp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN O2A1O1Ixp5_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.252 0.164 ;
        RECT 0.072 0.063 0.252 0.081 ;
        RECT 0.072 0.063 0.09 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.164 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.164 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.315 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.126 0.189 0.338 0.207 ;
      RECT 0.148 0.027 0.279 0.045 ;
      RECT 0.094 0.225 0.23 0.243 ;
  END
END O2A1O1Ixp5_ASAP7_75t_L

MACRO OA211x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211x2_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.09 0.144 ;
        RECT 0.018 0.07 0.036 0.2 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.164 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.296 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.286 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.252 0.243 ;
      RECT 0.234 0.189 0.252 0.243 ;
      RECT 0.234 0.189 0.306 0.207 ;
      RECT 0.288 0.063 0.306 0.207 ;
      RECT 0.099 0.063 0.306 0.081 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END OA211x2_ASAP7_75t_L

MACRO OA21x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21x2_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.07 0.036 0.236 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.153 0.239 0.171 ;
        RECT 0.18 0.106 0.198 0.171 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.225 0.36 0.243 ;
        RECT 0.342 0.027 0.36 0.243 ;
        RECT 0.256 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.148 0.225 0.224 0.243 ;
      RECT 0.206 0.189 0.224 0.243 ;
      RECT 0.206 0.189 0.306 0.207 ;
      RECT 0.288 0.063 0.306 0.207 ;
      RECT 0.099 0.063 0.306 0.081 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END OA21x2_ASAP7_75t_L

MACRO OA221x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221x2_ASAP7_75t_L 0 0 ;
  SIZE 0.864 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.215 0.189 0.252 0.207 ;
        RECT 0.234 0.099 0.252 0.207 ;
        RECT 0.215 0.099 0.252 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.189 0.379 0.207 ;
        RECT 0.342 0.099 0.379 0.117 ;
        RECT 0.342 0.099 0.36 0.207 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.593 0.189 0.63 0.207 ;
        RECT 0.612 0.099 0.63 0.207 ;
        RECT 0.593 0.099 0.63 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 0.189 0.522 0.207 ;
        RECT 0.504 0.099 0.522 0.207 ;
        RECT 0.485 0.099 0.522 0.117 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.189 0.757 0.207 ;
        RECT 0.72 0.099 0.757 0.117 ;
        RECT 0.72 0.099 0.738 0.207 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.864 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.122 0.045 ;
        RECT 0.018 0.225 0.117 0.243 ;
        RECT 0.099 0.189 0.117 0.243 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.144 0.225 0.846 0.243 ;
      RECT 0.828 0.063 0.846 0.243 ;
      RECT 0.144 0.126 0.162 0.243 ;
      RECT 0.121 0.126 0.162 0.144 ;
      RECT 0.741 0.063 0.846 0.081 ;
      RECT 0.472 0.027 0.824 0.045 ;
      RECT 0.202 0.063 0.668 0.081 ;
  END
END OA221x2_ASAP7_75t_L

MACRO OA222x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222x2_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.2 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.531 0.225 0.63 0.243 ;
        RECT 0.612 0.027 0.63 0.243 ;
        RECT 0.526 0.027 0.63 0.045 ;
        RECT 0.531 0.189 0.549 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.009 0.225 0.504 0.243 ;
      RECT 0.486 0.126 0.504 0.243 ;
      RECT 0.009 0.063 0.027 0.243 ;
      RECT 0.486 0.126 0.554 0.144 ;
      RECT 0.009 0.063 0.122 0.081 ;
      RECT 0.202 0.063 0.36 0.081 ;
      RECT 0.342 0.027 0.36 0.081 ;
      RECT 0.342 0.027 0.468 0.045 ;
      RECT 0.04 0.027 0.284 0.045 ;
  END
END OA222x2_ASAP7_75t_L

MACRO OA22x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22x2_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.236 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.063 0.414 0.2 ;
        RECT 0.367 0.063 0.414 0.081 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.071 0.225 0.122 0.243 ;
        RECT 0.071 0.027 0.122 0.045 ;
        RECT 0.071 0.027 0.091 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.225 0.392 0.243 ;
      RECT 0.18 0.063 0.198 0.243 ;
      RECT 0.137 0.126 0.198 0.144 ;
      RECT 0.18 0.063 0.333 0.081 ;
      RECT 0.256 0.027 0.5 0.045 ;
  END
END OA22x2_ASAP7_75t_L

MACRO OA31x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31x2_ASAP7_75t_L 0 0 ;
  SIZE 0.81 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.053 0.189 0.09 0.207 ;
        RECT 0.072 0.099 0.09 0.207 ;
        RECT 0.053 0.099 0.09 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.126 0.203 0.144 ;
        RECT 0.126 0.189 0.163 0.207 ;
        RECT 0.126 0.106 0.144 0.207 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.126 0.414 0.144 ;
        RECT 0.342 0.063 0.36 0.164 ;
        RECT 0.323 0.063 0.36 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 0.153 0.522 0.171 ;
        RECT 0.504 0.106 0.522 0.171 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.81 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.693 0.225 0.792 0.243 ;
        RECT 0.774 0.027 0.792 0.243 ;
        RECT 0.693 0.027 0.792 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.369 0.189 0.576 0.207 ;
      RECT 0.558 0.063 0.576 0.207 ;
      RECT 0.558 0.126 0.667 0.144 ;
      RECT 0.418 0.063 0.576 0.081 ;
      RECT 0.317 0.225 0.446 0.243 ;
      RECT 0.317 0.189 0.335 0.243 ;
      RECT 0.202 0.189 0.335 0.207 ;
      RECT 0.094 0.027 0.5 0.045 ;
      RECT 0.04 0.063 0.284 0.081 ;
      RECT 0.04 0.225 0.284 0.243 ;
  END
END OA31x2_ASAP7_75t_L

MACRO OA331x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA331x1_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.166 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.106 0.468 0.2 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.225 0.522 0.243 ;
      RECT 0.504 0.063 0.522 0.243 ;
      RECT 0.099 0.186 0.117 0.243 ;
      RECT 0.072 0.186 0.117 0.204 ;
      RECT 0.072 0.115 0.09 0.204 ;
      RECT 0.471 0.063 0.522 0.081 ;
      RECT 0.234 0.063 0.393 0.081 ;
      RECT 0.234 0.027 0.252 0.081 ;
      RECT 0.148 0.027 0.252 0.045 ;
      RECT 0.308 0.027 0.447 0.045 ;
  END
END OA331x1_ASAP7_75t_L

MACRO OA331x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA331x2_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.166 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.106 0.468 0.2 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.106 0.522 0.2 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.225 0.122 0.243 ;
        RECT 0.045 0.027 0.122 0.045 ;
        RECT 0.045 0.027 0.063 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.153 0.225 0.576 0.243 ;
      RECT 0.558 0.063 0.576 0.243 ;
      RECT 0.153 0.186 0.171 0.243 ;
      RECT 0.126 0.186 0.171 0.204 ;
      RECT 0.126 0.115 0.144 0.204 ;
      RECT 0.525 0.063 0.576 0.081 ;
      RECT 0.288 0.063 0.447 0.081 ;
      RECT 0.288 0.027 0.306 0.081 ;
      RECT 0.202 0.027 0.306 0.045 ;
      RECT 0.362 0.027 0.501 0.045 ;
  END
END OA331x2_ASAP7_75t_L

MACRO OA332x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA332x1_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.106 0.522 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.106 0.468 0.2 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.094 0.243 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.126 0.225 0.576 0.243 ;
      RECT 0.558 0.063 0.576 0.243 ;
      RECT 0.126 0.189 0.144 0.243 ;
      RECT 0.072 0.189 0.144 0.207 ;
      RECT 0.072 0.119 0.09 0.207 ;
      RECT 0.471 0.063 0.576 0.081 ;
      RECT 0.234 0.063 0.393 0.081 ;
      RECT 0.234 0.027 0.252 0.081 ;
      RECT 0.146 0.027 0.252 0.045 ;
      RECT 0.308 0.027 0.556 0.045 ;
  END
END OA332x1_ASAP7_75t_L

MACRO OA332x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA332x2_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.106 0.468 0.2 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.106 0.576 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.106 0.522 0.2 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.137 0.243 ;
        RECT 0.018 0.027 0.122 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.225 0.63 0.243 ;
      RECT 0.612 0.063 0.63 0.243 ;
      RECT 0.18 0.189 0.198 0.243 ;
      RECT 0.126 0.189 0.198 0.207 ;
      RECT 0.126 0.119 0.144 0.207 ;
      RECT 0.525 0.063 0.63 0.081 ;
      RECT 0.288 0.063 0.447 0.081 ;
      RECT 0.288 0.027 0.306 0.081 ;
      RECT 0.2 0.027 0.306 0.045 ;
      RECT 0.362 0.027 0.61 0.045 ;
  END
END OA332x2_ASAP7_75t_L

MACRO OA333x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA333x1_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.106 0.576 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.106 0.522 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.106 0.468 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.164 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.225 0.63 0.243 ;
      RECT 0.612 0.063 0.63 0.243 ;
      RECT 0.099 0.186 0.117 0.243 ;
      RECT 0.072 0.186 0.117 0.204 ;
      RECT 0.072 0.115 0.09 0.204 ;
      RECT 0.467 0.063 0.63 0.081 ;
      RECT 0.232 0.063 0.394 0.081 ;
      RECT 0.232 0.027 0.25 0.081 ;
      RECT 0.147 0.027 0.25 0.045 ;
      RECT 0.309 0.027 0.569 0.045 ;
  END
END OA333x1_ASAP7_75t_L

MACRO OA333x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA333x2_ASAP7_75t_L 0 0 ;
  SIZE 0.702 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.106 0.63 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.106 0.576 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.106 0.522 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.106 0.468 0.2 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.164 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.702 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.225 0.122 0.243 ;
        RECT 0.072 0.027 0.122 0.045 ;
        RECT 0.072 0.027 0.09 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.153 0.225 0.684 0.243 ;
      RECT 0.666 0.063 0.684 0.243 ;
      RECT 0.153 0.186 0.171 0.243 ;
      RECT 0.126 0.186 0.171 0.204 ;
      RECT 0.126 0.115 0.144 0.204 ;
      RECT 0.521 0.063 0.684 0.081 ;
      RECT 0.286 0.063 0.448 0.081 ;
      RECT 0.286 0.027 0.304 0.081 ;
      RECT 0.201 0.027 0.304 0.045 ;
      RECT 0.363 0.027 0.623 0.045 ;
  END
END OA333x2_ASAP7_75t_L

MACRO OA33x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA33x2_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.106 0.468 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.122 0.045 ;
        RECT 0.018 0.225 0.117 0.243 ;
        RECT 0.099 0.189 0.117 0.243 ;
        RECT 0.062 0.189 0.117 0.207 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.144 0.225 0.522 0.243 ;
      RECT 0.504 0.063 0.522 0.243 ;
      RECT 0.144 0.126 0.162 0.243 ;
      RECT 0.121 0.126 0.162 0.144 ;
      RECT 0.364 0.063 0.522 0.081 ;
      RECT 0.202 0.027 0.446 0.045 ;
  END
END OA33x2_ASAP7_75t_L

MACRO OAI211xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.09 0.144 ;
        RECT 0.018 0.07 0.036 0.2 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.04 0.225 0.306 0.243 ;
        RECT 0.288 0.063 0.306 0.243 ;
        RECT 0.099 0.063 0.306 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END OAI211xp5_ASAP7_75t_L

MACRO OAI21x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21x1_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.189 0.306 0.207 ;
        RECT 0.288 0.106 0.306 0.207 ;
        RECT 0.126 0.106 0.144 0.207 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.19 0.127 0.256 0.145 ;
        RECT 0.19 0.099 0.227 0.171 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.063 0.36 0.154 ;
        RECT 0.072 0.063 0.36 0.081 ;
        RECT 0.072 0.063 0.09 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.369 0.027 0.414 0.045 ;
        RECT 0.018 0.027 0.063 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.027 0.333 0.045 ;
  END
END OAI21x1_ASAP7_75t_L

MACRO OAI21xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.27 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.07 0.036 0.236 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.203 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.27 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.225 0.252 0.243 ;
        RECT 0.234 0.063 0.252 0.243 ;
        RECT 0.099 0.063 0.252 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END OAI21xp33_ASAP7_75t_L

MACRO OAI21xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.27 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.07 0.036 0.236 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.203 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.171 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.27 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.225 0.252 0.243 ;
        RECT 0.234 0.063 0.252 0.243 ;
        RECT 0.099 0.063 0.252 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END OAI21xp5_ASAP7_75t_L

MACRO OAI221xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.236 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.23 0.243 ;
        RECT 0.018 0.063 0.123 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.201 0.063 0.339 0.081 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END OAI221xp5_ASAP7_75t_L

MACRO OAI222xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.07 0.414 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.07 0.468 0.2 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.522 0.243 ;
        RECT 0.504 0.055 0.522 0.243 ;
        RECT 0.018 0.063 0.122 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.063 0.36 0.081 ;
      RECT 0.342 0.027 0.36 0.081 ;
      RECT 0.342 0.027 0.468 0.045 ;
      RECT 0.04 0.027 0.284 0.045 ;
  END
END OAI222xp33_ASAP7_75t_L

MACRO OAI22x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22x1_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.153 0.379 0.171 ;
        RECT 0.342 0.099 0.379 0.117 ;
        RECT 0.342 0.099 0.36 0.171 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.189 0.468 0.207 ;
        RECT 0.45 0.099 0.468 0.207 ;
        RECT 0.431 0.099 0.468 0.117 ;
        RECT 0.288 0.118 0.306 0.207 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.161 0.153 0.198 0.171 ;
        RECT 0.18 0.063 0.198 0.171 ;
        RECT 0.161 0.063 0.198 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.189 0.252 0.207 ;
        RECT 0.234 0.116 0.252 0.207 ;
        RECT 0.072 0.063 0.109 0.081 ;
        RECT 0.072 0.063 0.09 0.207 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.038 0.225 0.522 0.243 ;
        RECT 0.504 0.063 0.522 0.243 ;
        RECT 0.309 0.063 0.522 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.5 0.045 ;
  END
END OAI22x1_ASAP7_75t_L

MACRO OAI22xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.225 0.275 0.243 ;
        RECT 0.234 0.07 0.252 0.243 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.176 0.243 ;
        RECT 0.018 0.063 0.117 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.284 0.045 ;
  END
END OAI22xp33_ASAP7_75t_L

MACRO OAI22xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.225 0.275 0.243 ;
        RECT 0.234 0.07 0.252 0.243 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.063 0.198 0.164 ;
        RECT 0.151 0.063 0.198 0.081 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.176 0.243 ;
        RECT 0.018 0.063 0.117 0.081 ;
        RECT 0.018 0.063 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.284 0.045 ;
  END
END OAI22xp5_ASAP7_75t_L

MACRO OAI311xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI311xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.236 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.2 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.2 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.198 0.225 0.36 0.243 ;
        RECT 0.342 0.027 0.36 0.243 ;
        RECT 0.31 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.027 0.234 0.045 ;
  END
END OAI311xp33_ASAP7_75t_L

MACRO OAI31xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.236 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.236 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.201 0.225 0.306 0.243 ;
        RECT 0.288 0.063 0.306 0.243 ;
        RECT 0.256 0.063 0.306 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.093 0.027 0.23 0.045 ;
  END
END OAI31xp33_ASAP7_75t_L

MACRO OAI31xp67_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31xp67_ASAP7_75t_L 0 0 ;
  SIZE 0.702 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.666 0.126 0.684 0.198 ;
        RECT 0.553 0.126 0.684 0.144 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.126 0.419 0.144 ;
        RECT 0.288 0.126 0.306 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.07 0.036 0.236 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.126 0.203 0.144 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.702 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.063 0.663 0.081 ;
        RECT 0.202 0.189 0.252 0.207 ;
        RECT 0.234 0.063 0.252 0.207 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.526 0.225 0.663 0.243 ;
      RECT 0.364 0.189 0.608 0.207 ;
      RECT 0.04 0.027 0.554 0.045 ;
      RECT 0.094 0.225 0.446 0.243 ;
  END
END OAI31xp67_ASAP7_75t_L

MACRO OAI321xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI321xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.236 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.095 0.144 ;
        RECT 0.018 0.034 0.036 0.236 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.198 0.225 0.414 0.243 ;
        RECT 0.396 0.063 0.414 0.243 ;
        RECT 0.31 0.063 0.414 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.256 0.027 0.396 0.045 ;
      RECT 0.094 0.063 0.23 0.081 ;
  END
END OAI321xp33_ASAP7_75t_L

MACRO OAI322xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI322xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.105 0.306 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.236 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.105 0.36 0.2 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.147 0.225 0.468 0.243 ;
        RECT 0.45 0.063 0.468 0.243 ;
        RECT 0.364 0.063 0.468 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.027 0.45 0.045 ;
      RECT 0.039 0.063 0.284 0.081 ;
  END
END OAI322xp33_ASAP7_75t_L

MACRO OAI32xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.063 0.222 0.081 ;
        RECT 0.18 0.063 0.198 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.04 0.225 0.36 0.243 ;
        RECT 0.342 0.063 0.36 0.243 ;
        RECT 0.256 0.063 0.36 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.027 0.338 0.045 ;
  END
END OAI32xp33_ASAP7_75t_L

MACRO OAI331xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI331xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.236 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.236 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.201 0.225 0.468 0.243 ;
        RECT 0.45 0.063 0.468 0.243 ;
        RECT 0.417 0.063 0.468 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.254 0.027 0.393 0.045 ;
      RECT 0.092 0.063 0.339 0.081 ;
  END
END OAI331xp33_ASAP7_75t_L

MACRO OAI332xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI332xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.54 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.236 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.236 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.106 0.468 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.54 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.201 0.225 0.522 0.243 ;
        RECT 0.504 0.063 0.522 0.243 ;
        RECT 0.417 0.063 0.522 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.254 0.027 0.502 0.045 ;
      RECT 0.092 0.063 0.339 0.081 ;
  END
END OAI332xp33_ASAP7_75t_L

MACRO OAI333xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI333xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.106 0.522 0.2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.106 0.468 0.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.236 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.106 0.09 0.236 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.201 0.225 0.576 0.243 ;
        RECT 0.558 0.063 0.576 0.243 ;
        RECT 0.413 0.063 0.576 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.254 0.027 0.515 0.045 ;
      RECT 0.094 0.063 0.34 0.081 ;
  END
END OAI333xp33_ASAP7_75t_L

MACRO OAI33xp33_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33xp33_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.236 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.236 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.106 0.252 0.2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.2 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.106 0.36 0.2 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.201 0.225 0.414 0.243 ;
        RECT 0.396 0.063 0.414 0.243 ;
        RECT 0.256 0.063 0.414 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.092 0.027 0.338 0.045 ;
  END
END OAI33xp33_ASAP7_75t_L

MACRO OR2x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x2_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.077 0.144 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.225 0.306 0.243 ;
        RECT 0.288 0.027 0.306 0.243 ;
        RECT 0.207 0.027 0.306 0.045 ;
        RECT 0.207 0.184 0.225 0.243 ;
        RECT 0.207 0.027 0.225 0.086 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.186 0.243 ;
      RECT 0.168 0.027 0.186 0.243 ;
      RECT 0.168 0.126 0.227 0.144 ;
      RECT 0.094 0.027 0.186 0.045 ;
  END
END OR2x2_ASAP7_75t_L

MACRO OR2x4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x4_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.126 0.077 0.144 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.207 0.027 0.414 0.045 ;
        RECT 0.315 0.184 0.333 0.243 ;
        RECT 0.315 0.027 0.333 0.086 ;
        RECT 0.207 0.184 0.225 0.243 ;
        RECT 0.207 0.027 0.225 0.086 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.187 0.243 ;
      RECT 0.169 0.027 0.187 0.243 ;
      RECT 0.169 0.126 0.227 0.144 ;
      RECT 0.094 0.027 0.187 0.045 ;
  END
END OR2x4_ASAP7_75t_L

MACRO OR2x6_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x6_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.063 0.144 0.122 ;
        RECT 0.018 0.063 0.144 0.081 ;
        RECT 0.018 0.063 0.036 0.236 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.153 0.252 0.171 ;
        RECT 0.234 0.121 0.252 0.171 ;
        RECT 0.072 0.106 0.09 0.236 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.225 0.63 0.243 ;
        RECT 0.612 0.027 0.63 0.243 ;
        RECT 0.31 0.027 0.63 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.148 0.189 0.306 0.207 ;
      RECT 0.288 0.07 0.306 0.207 ;
      RECT 0.234 0.07 0.306 0.088 ;
      RECT 0.234 0.027 0.252 0.088 ;
      RECT 0.094 0.027 0.252 0.045 ;
  END
END OR2x6_ASAP7_75t_L

MACRO OR3x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x1_ASAP7_75t_L 0 0 ;
  SIZE 0.324 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.324 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.183 0.306 0.201 ;
        RECT 0.288 0.076 0.306 0.201 ;
        RECT 0.261 0.076 0.306 0.094 ;
        RECT 0.261 0.183 0.279 0.235 ;
        RECT 0.261 0.034 0.279 0.094 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.234 0.243 ;
      RECT 0.216 0.027 0.234 0.243 ;
      RECT 0.216 0.126 0.262 0.144 ;
      RECT 0.04 0.027 0.234 0.045 ;
  END
END OR3x1_ASAP7_75t_L

MACRO OR3x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x2_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.225 0.36 0.243 ;
        RECT 0.342 0.027 0.36 0.243 ;
        RECT 0.261 0.027 0.36 0.045 ;
        RECT 0.261 0.184 0.279 0.243 ;
        RECT 0.261 0.027 0.279 0.086 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.24 0.243 ;
      RECT 0.222 0.027 0.24 0.243 ;
      RECT 0.222 0.126 0.284 0.144 ;
      RECT 0.04 0.027 0.24 0.045 ;
  END
END OR3x2_ASAP7_75t_L

MACRO OR3x4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x4_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.2 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.261 0.027 0.468 0.045 ;
        RECT 0.369 0.184 0.387 0.243 ;
        RECT 0.369 0.027 0.387 0.086 ;
        RECT 0.261 0.184 0.279 0.243 ;
        RECT 0.261 0.027 0.279 0.086 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.225 0.241 0.243 ;
      RECT 0.223 0.027 0.241 0.243 ;
      RECT 0.223 0.126 0.284 0.144 ;
      RECT 0.04 0.027 0.241 0.045 ;
  END
END OR3x4_ASAP7_75t_L

MACRO OR4x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4x1_ASAP7_75t_L 0 0 ;
  SIZE 0.378 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.236 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.236 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.106 0.144 0.236 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.378 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.31 0.225 0.36 0.243 ;
      RECT 0.342 0.027 0.36 0.243 ;
      RECT 0.072 0.066 0.09 0.152 ;
      RECT 0.072 0.066 0.117 0.084 ;
      RECT 0.099 0.027 0.117 0.084 ;
      RECT 0.099 0.027 0.36 0.045 ;
  END
END OR4x1_ASAP7_75t_L

MACRO OR4x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4x2_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.07 0.36 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.07 0.306 0.236 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.236 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.106 0.198 0.236 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.122 0.243 ;
        RECT 0.018 0.027 0.122 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.225 0.414 0.243 ;
      RECT 0.396 0.027 0.414 0.243 ;
      RECT 0.099 0.063 0.117 0.149 ;
      RECT 0.099 0.063 0.171 0.081 ;
      RECT 0.153 0.027 0.171 0.081 ;
      RECT 0.153 0.027 0.414 0.045 ;
  END
END OR4x2_ASAP7_75t_L

MACRO OR5x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5x1_ASAP7_75t_L 0 0 ;
  SIZE 0.432 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.236 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.236 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.236 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.236 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.432 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.35 0.225 0.414 0.243 ;
        RECT 0.396 0.027 0.414 0.243 ;
        RECT 0.349 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.225 0.07 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.342 0.063 0.36 0.154 ;
      RECT 0.288 0.063 0.36 0.081 ;
      RECT 0.288 0.027 0.306 0.081 ;
      RECT 0.018 0.027 0.306 0.045 ;
  END
END OR5x1_ASAP7_75t_L

MACRO OR5x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5x2_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.07 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.236 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.236 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.07 0.252 0.236 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.106 0.306 0.236 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.343 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.225 0.07 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.342 0.063 0.36 0.154 ;
      RECT 0.288 0.063 0.36 0.081 ;
      RECT 0.288 0.027 0.306 0.081 ;
      RECT 0.018 0.027 0.306 0.045 ;
  END
END OR5x2_ASAP7_75t_L

MACRO SDFHx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFHx1_ASAP7_75t_L 0 0 ;
  SIZE 1.35 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.282 0.225 1.332 0.243 ;
        RECT 1.314 0.027 1.332 0.243 ;
        RECT 1.282 0.027 1.332 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.35 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.211 0.036 1.229 0.054 ;
      LAYER M1 ;
        RECT 1.206 0.027 1.25 0.045 ;
        RECT 1.206 0.027 1.224 0.2 ;
        RECT 0.216 0.126 0.311 0.144 ;
        RECT 0.216 0.027 0.258 0.045 ;
        RECT 0.216 0.027 0.234 0.144 ;
      LAYER V1 ;
        RECT 0.216 0.036 0.234 0.054 ;
        RECT 1.206 0.036 1.224 0.054 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.467 0.108 0.59 0.126 ;
      LAYER M1 ;
        RECT 0.485 0.189 0.522 0.207 ;
        RECT 0.504 0.106 0.522 0.207 ;
        RECT 0.461 0.126 0.522 0.144 ;
      LAYER V1 ;
        RECT 0.504 0.108 0.522 0.126 ;
    END
  END SI
  OBS
    LAYER M1 ;
      RECT 1.152 0.225 1.202 0.243 ;
      RECT 1.152 0.034 1.17 0.243 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.342 0.063 0.36 0.164 ;
      RECT 0.342 0.063 0.379 0.081 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.26 0.09 1.278 0.2 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.283 0.162 ;
      RECT 0.337 0.072 1.175 0.09 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.175 0.18 0.743 0.198 ;
    LAYER V1 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.152 0.072 1.17 0.09 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.342 0.072 0.36 0.09 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
  END
END SDFHx1_ASAP7_75t_L

MACRO SDFHx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFHx2_ASAP7_75t_L 0 0 ;
  SIZE 1.404 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.081 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.099 0.433 0.117 ;
        RECT 0.396 0.099 0.414 0.164 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.282 0.225 1.386 0.243 ;
        RECT 1.368 0.027 1.386 0.243 ;
        RECT 1.282 0.027 1.386 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.211 0.036 1.229 0.054 ;
      LAYER M1 ;
        RECT 1.206 0.027 1.25 0.045 ;
        RECT 1.206 0.027 1.224 0.2 ;
        RECT 0.216 0.126 0.311 0.144 ;
        RECT 0.216 0.027 0.258 0.045 ;
        RECT 0.216 0.027 0.234 0.144 ;
      LAYER V1 ;
        RECT 0.216 0.036 0.234 0.054 ;
        RECT 1.206 0.036 1.224 0.054 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 0.189 0.522 0.207 ;
        RECT 0.504 0.106 0.522 0.207 ;
        RECT 0.461 0.126 0.522 0.144 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.404 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.152 0.225 1.202 0.243 ;
      RECT 1.152 0.034 1.17 0.243 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.792 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.342 0.063 0.36 0.164 ;
      RECT 0.342 0.063 0.379 0.081 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 1.26 0.09 1.278 0.2 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.283 0.162 ;
      RECT 0.337 0.072 1.175 0.09 ;
      RECT 0.019 0.144 0.9 0.162 ;
      RECT 0.175 0.18 0.743 0.198 ;
    LAYER V1 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.152 0.072 1.17 0.09 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.342 0.072 0.36 0.09 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END SDFHx2_ASAP7_75t_L

MACRO SDFHx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFHx3_ASAP7_75t_L 0 0 ;
  SIZE 1.458 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.081 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.099 0.433 0.117 ;
        RECT 0.396 0.099 0.414 0.164 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.282 0.225 1.44 0.243 ;
        RECT 1.422 0.027 1.44 0.243 ;
        RECT 1.282 0.027 1.44 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.211 0.036 1.229 0.054 ;
      LAYER M1 ;
        RECT 1.206 0.027 1.25 0.045 ;
        RECT 1.206 0.027 1.224 0.2 ;
        RECT 0.216 0.126 0.311 0.144 ;
        RECT 0.216 0.027 0.258 0.045 ;
        RECT 0.216 0.027 0.234 0.144 ;
      LAYER V1 ;
        RECT 0.216 0.036 0.234 0.054 ;
        RECT 1.206 0.036 1.224 0.054 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 0.189 0.522 0.207 ;
        RECT 0.504 0.106 0.522 0.207 ;
        RECT 0.461 0.126 0.522 0.144 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.458 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.458 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.152 0.225 1.202 0.243 ;
      RECT 1.152 0.034 1.17 0.243 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.792 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.342 0.063 0.36 0.164 ;
      RECT 0.342 0.063 0.379 0.081 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 1.26 0.09 1.278 0.2 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.283 0.162 ;
      RECT 0.337 0.072 1.175 0.09 ;
      RECT 0.019 0.144 0.9 0.162 ;
      RECT 0.175 0.18 0.743 0.198 ;
    LAYER V1 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.152 0.072 1.17 0.09 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.342 0.072 0.36 0.09 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END SDFHx3_ASAP7_75t_L

MACRO SDFHx4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFHx4_ASAP7_75t_L 0 0 ;
  SIZE 1.674 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.063 0.109 0.081 ;
        RECT 0.072 0.063 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.099 0.468 0.164 ;
        RECT 0.378 0.225 0.459 0.243 ;
        RECT 0.378 0.099 0.468 0.117 ;
        RECT 0.378 0.099 0.396 0.243 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.444 0.225 1.656 0.243 ;
        RECT 1.637 0.027 1.656 0.243 ;
        RECT 1.444 0.027 1.656 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.229 0.072 0.581 0.09 ;
      LAYER M1 ;
        RECT 0.558 0.063 0.599 0.081 ;
        RECT 0.558 0.063 0.576 0.164 ;
        RECT 0.234 0.126 0.289 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
      LAYER V1 ;
        RECT 0.234 0.072 0.252 0.09 ;
        RECT 0.558 0.072 0.576 0.09 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.693 0.027 0.767 0.045 ;
        RECT 0.639 0.063 0.711 0.081 ;
        RECT 0.693 0.027 0.711 0.081 ;
        RECT 0.612 0.106 0.657 0.124 ;
        RECT 0.639 0.063 0.657 0.124 ;
        RECT 0.612 0.106 0.63 0.164 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.674 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.674 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.059 0.225 1.386 0.243 ;
      RECT 1.368 0.027 1.386 0.243 ;
      RECT 1.368 0.126 1.447 0.144 ;
      RECT 1.242 0.126 1.283 0.144 ;
      RECT 1.242 0.027 1.26 0.144 ;
      RECT 1.113 0.027 1.386 0.045 ;
      RECT 1.206 0.182 1.332 0.2 ;
      RECT 1.314 0.081 1.332 0.2 ;
      RECT 1.206 0.106 1.224 0.2 ;
      RECT 1.287 0.081 1.332 0.099 ;
      RECT 0.882 0.063 0.9 0.164 ;
      RECT 0.882 0.063 0.981 0.081 ;
      RECT 0.801 0.225 0.954 0.243 ;
      RECT 0.936 0.106 0.954 0.243 ;
      RECT 0.801 0.189 0.819 0.243 ;
      RECT 0.738 0.189 0.819 0.207 ;
      RECT 0.738 0.07 0.756 0.207 ;
      RECT 0.31 0.225 0.36 0.243 ;
      RECT 0.342 0.027 0.36 0.243 ;
      RECT 0.504 0.063 0.522 0.164 ;
      RECT 0.342 0.063 0.522 0.081 ;
      RECT 0.31 0.027 0.36 0.045 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.126 0.027 0.198 0.045 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.09 0.045 ;
      RECT 1.152 0.106 1.17 0.2 ;
      RECT 1.098 0.07 1.116 0.164 ;
      RECT 1.044 0.106 1.062 0.2 ;
      RECT 0.828 0.07 0.846 0.167 ;
      RECT 0.774 0.07 0.792 0.164 ;
      RECT 0.58 0.225 0.77 0.243 ;
      RECT 0.684 0.121 0.702 0.167 ;
      RECT 0.418 0.027 0.662 0.045 ;
      RECT 0.423 0.189 0.662 0.207 ;
      RECT 0.126 0.106 0.144 0.2 ;
    LAYER M2 ;
      RECT 0.019 0.144 1.175 0.162 ;
      RECT 0.175 0.108 1.121 0.126 ;
    LAYER V1 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.098 0.108 1.116 0.126 ;
      RECT 1.044 0.144 1.062 0.162 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.774 0.108 0.792 0.126 ;
      RECT 0.684 0.144 0.702 0.162 ;
      RECT 0.18 0.108 0.198 0.126 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.024 0.144 0.042 0.162 ;
  END
END SDFHx4_ASAP7_75t_L

MACRO SDFLx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx1_ASAP7_75t_L 0 0 ;
  SIZE 1.35 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.081 0.09 0.164 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.099 0.433 0.117 ;
        RECT 0.396 0.099 0.414 0.164 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.282 0.225 1.332 0.243 ;
        RECT 1.314 0.027 1.332 0.243 ;
        RECT 1.282 0.027 1.332 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.211 0.036 1.229 0.054 ;
      LAYER M1 ;
        RECT 1.206 0.027 1.25 0.045 ;
        RECT 1.206 0.027 1.224 0.2 ;
        RECT 0.216 0.126 0.311 0.144 ;
        RECT 0.216 0.027 0.258 0.045 ;
        RECT 0.216 0.027 0.234 0.144 ;
      LAYER V1 ;
        RECT 0.216 0.036 0.234 0.054 ;
        RECT 1.206 0.036 1.224 0.054 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 0.189 0.522 0.207 ;
        RECT 0.504 0.106 0.522 0.207 ;
        RECT 0.461 0.126 0.522 0.144 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.35 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.152 0.225 1.202 0.243 ;
      RECT 1.152 0.034 1.17 0.243 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.342 0.063 0.36 0.164 ;
      RECT 0.342 0.063 0.379 0.081 ;
      RECT 0.126 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.107 0.189 0.144 0.207 ;
      RECT 0.126 0.121 0.144 0.207 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 1.26 0.09 1.278 0.2 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.309 0.189 0.447 0.207 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.283 0.162 ;
      RECT 0.337 0.072 1.175 0.09 ;
      RECT 0.175 0.144 0.9 0.162 ;
      RECT 0.019 0.18 0.743 0.198 ;
    LAYER V1 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.152 0.072 1.17 0.09 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.342 0.072 0.36 0.09 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.126 0.18 0.144 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END SDFLx1_ASAP7_75t_L

MACRO SDFLx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx2_ASAP7_75t_L 0 0 ;
  SIZE 1.404 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.081 0.09 0.164 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.099 0.433 0.117 ;
        RECT 0.396 0.099 0.414 0.164 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.282 0.225 1.386 0.243 ;
        RECT 1.368 0.027 1.386 0.243 ;
        RECT 1.282 0.027 1.386 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.211 0.036 1.229 0.054 ;
      LAYER M1 ;
        RECT 1.206 0.027 1.25 0.045 ;
        RECT 1.206 0.027 1.224 0.2 ;
        RECT 0.216 0.126 0.311 0.144 ;
        RECT 0.216 0.027 0.258 0.045 ;
        RECT 0.216 0.027 0.234 0.144 ;
      LAYER V1 ;
        RECT 0.216 0.036 0.234 0.054 ;
        RECT 1.206 0.036 1.224 0.054 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 0.189 0.522 0.207 ;
        RECT 0.504 0.106 0.522 0.207 ;
        RECT 0.461 0.126 0.522 0.144 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.404 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.152 0.225 1.202 0.243 ;
      RECT 1.152 0.034 1.17 0.243 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.792 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.342 0.063 0.36 0.164 ;
      RECT 0.342 0.063 0.379 0.081 ;
      RECT 0.126 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.107 0.189 0.144 0.207 ;
      RECT 0.126 0.121 0.144 0.207 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 1.26 0.09 1.278 0.2 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.309 0.189 0.447 0.207 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.283 0.162 ;
      RECT 0.337 0.072 1.175 0.09 ;
      RECT 0.175 0.144 0.9 0.162 ;
      RECT 0.019 0.18 0.743 0.198 ;
    LAYER V1 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.152 0.072 1.17 0.09 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.342 0.072 0.36 0.09 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.126 0.18 0.144 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END SDFLx2_ASAP7_75t_L

MACRO SDFLx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx3_ASAP7_75t_L 0 0 ;
  SIZE 1.458 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.081 0.09 0.164 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.099 0.433 0.117 ;
        RECT 0.396 0.099 0.414 0.164 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.282 0.225 1.44 0.243 ;
        RECT 1.422 0.027 1.44 0.243 ;
        RECT 1.282 0.027 1.44 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.211 0.036 1.229 0.054 ;
      LAYER M1 ;
        RECT 1.206 0.027 1.25 0.045 ;
        RECT 1.206 0.027 1.224 0.2 ;
        RECT 0.216 0.126 0.311 0.144 ;
        RECT 0.216 0.027 0.258 0.045 ;
        RECT 0.216 0.027 0.234 0.144 ;
      LAYER V1 ;
        RECT 0.216 0.036 0.234 0.054 ;
        RECT 1.206 0.036 1.224 0.054 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 0.189 0.522 0.207 ;
        RECT 0.504 0.106 0.522 0.207 ;
        RECT 0.461 0.126 0.522 0.144 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.458 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.458 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.152 0.225 1.202 0.243 ;
      RECT 1.152 0.034 1.17 0.243 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.792 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.342 0.063 0.36 0.164 ;
      RECT 0.342 0.063 0.379 0.081 ;
      RECT 0.126 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.107 0.189 0.144 0.207 ;
      RECT 0.126 0.121 0.144 0.207 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.18 0.047 0.198 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 1.26 0.09 1.278 0.2 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.309 0.189 0.447 0.207 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.283 0.162 ;
      RECT 0.337 0.072 1.175 0.09 ;
      RECT 0.175 0.144 0.9 0.162 ;
      RECT 0.019 0.18 0.743 0.198 ;
    LAYER V1 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.152 0.072 1.17 0.09 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.342 0.072 0.36 0.09 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.126 0.18 0.144 0.198 ;
      RECT 0.024 0.18 0.042 0.198 ;
  END
END SDFLx3_ASAP7_75t_L

MACRO SDFLx4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx4_ASAP7_75t_L 0 0 ;
  SIZE 1.674 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.063 0.109 0.081 ;
        RECT 0.072 0.063 0.09 0.2 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.099 0.468 0.164 ;
        RECT 0.378 0.225 0.459 0.243 ;
        RECT 0.378 0.099 0.468 0.117 ;
        RECT 0.378 0.099 0.396 0.243 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.444 0.225 1.656 0.243 ;
        RECT 1.637 0.027 1.656 0.243 ;
        RECT 1.444 0.027 1.656 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.229 0.072 0.581 0.09 ;
      LAYER M1 ;
        RECT 0.558 0.063 0.599 0.081 ;
        RECT 0.558 0.063 0.576 0.164 ;
        RECT 0.234 0.126 0.289 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
      LAYER V1 ;
        RECT 0.234 0.072 0.252 0.09 ;
        RECT 0.558 0.072 0.576 0.09 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.693 0.027 0.767 0.045 ;
        RECT 0.639 0.063 0.711 0.081 ;
        RECT 0.693 0.027 0.711 0.081 ;
        RECT 0.612 0.106 0.657 0.124 ;
        RECT 0.639 0.063 0.657 0.124 ;
        RECT 0.612 0.106 0.63 0.164 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.674 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.674 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.059 0.225 1.386 0.243 ;
      RECT 1.368 0.027 1.386 0.243 ;
      RECT 1.368 0.126 1.447 0.144 ;
      RECT 1.242 0.126 1.283 0.144 ;
      RECT 1.242 0.027 1.26 0.144 ;
      RECT 1.113 0.027 1.386 0.045 ;
      RECT 1.206 0.182 1.332 0.2 ;
      RECT 1.314 0.081 1.332 0.2 ;
      RECT 1.206 0.106 1.224 0.2 ;
      RECT 1.287 0.081 1.332 0.099 ;
      RECT 0.882 0.063 0.9 0.164 ;
      RECT 0.882 0.063 0.981 0.081 ;
      RECT 0.801 0.225 0.954 0.243 ;
      RECT 0.936 0.106 0.954 0.243 ;
      RECT 0.801 0.189 0.819 0.243 ;
      RECT 0.738 0.189 0.819 0.207 ;
      RECT 0.738 0.07 0.756 0.207 ;
      RECT 0.31 0.225 0.36 0.243 ;
      RECT 0.342 0.027 0.36 0.243 ;
      RECT 0.504 0.063 0.522 0.164 ;
      RECT 0.342 0.063 0.522 0.081 ;
      RECT 0.31 0.027 0.36 0.045 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.126 0.027 0.198 0.045 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.108 0.047 0.126 ;
      RECT 0.009 0.027 0.09 0.045 ;
      RECT 1.152 0.106 1.17 0.2 ;
      RECT 1.098 0.07 1.116 0.164 ;
      RECT 1.044 0.106 1.062 0.2 ;
      RECT 0.828 0.07 0.846 0.167 ;
      RECT 0.774 0.07 0.792 0.164 ;
      RECT 0.58 0.225 0.77 0.243 ;
      RECT 0.684 0.121 0.702 0.167 ;
      RECT 0.418 0.027 0.662 0.045 ;
      RECT 0.423 0.189 0.662 0.207 ;
      RECT 0.126 0.103 0.144 0.2 ;
    LAYER M2 ;
      RECT 0.175 0.144 1.175 0.162 ;
      RECT 0.019 0.108 1.121 0.126 ;
    LAYER V1 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.098 0.108 1.116 0.126 ;
      RECT 1.044 0.144 1.062 0.162 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.774 0.108 0.792 0.126 ;
      RECT 0.684 0.144 0.702 0.162 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.126 0.108 0.144 0.126 ;
      RECT 0.024 0.108 0.042 0.126 ;
  END
END SDFLx4_ASAP7_75t_L

MACRO TAPCELL_ASAP7_75t_L
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN TAPCELL_ASAP7_75t_L 0 0 ;
  SIZE 0.108 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.108 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.108 0.009 ;
    END
  END VSS
END TAPCELL_ASAP7_75t_L

MACRO TAPCELL_WITH_FILLER_ASAP7_75t_L
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN TAPCELL_WITH_FILLER_ASAP7_75t_L 0 0 ;
  SIZE 0.162 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.162 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
END TAPCELL_WITH_FILLER_ASAP7_75t_L

MACRO TIEHIx1_ASAP7_75t_L
  CLASS CORE TIEHIGH ;
  ORIGIN 0 0 ;
  FOREIGN TIEHIx1_ASAP7_75t_L 0 0 ;
  SIZE 0.162 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.225 0.144 0.243 ;
        RECT 0.126 0.07 0.144 0.243 ;
        RECT 0.067 0.07 0.144 0.088 ;
    END
  END H
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.162 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.018 0.128 0.095 0.146 ;
      RECT 0.018 0.027 0.036 0.146 ;
      RECT 0.018 0.027 0.068 0.045 ;
  END
END TIEHIx1_ASAP7_75t_L

MACRO TIELOx1_ASAP7_75t_L
  CLASS CORE TIELOW ;
  ORIGIN 0 0 ;
  FOREIGN TIELOx1_ASAP7_75t_L 0 0 ;
  SIZE 0.162 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN L
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.067 0.182 0.144 0.2 ;
        RECT 0.126 0.027 0.144 0.2 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END L
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.162 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.124 0.036 0.243 ;
      RECT 0.018 0.124 0.095 0.142 ;
  END
END TIELOx1_ASAP7_75t_L

MACRO XNOR2x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x1_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.298 0.072 0.527 0.09 ;
      LAYER M1 ;
        RECT 0.504 0.07 0.522 0.152 ;
        RECT 0.305 0.126 0.365 0.144 ;
        RECT 0.305 0.067 0.323 0.144 ;
        RECT 0.213 0.067 0.323 0.085 ;
        RECT 0.213 0.027 0.231 0.085 ;
        RECT 0.018 0.027 0.231 0.045 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.027 0.036 0.236 ;
      LAYER V1 ;
        RECT 0.305 0.072 0.323 0.09 ;
        RECT 0.504 0.072 0.522 0.09 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.225 0.612 0.243 ;
        RECT 0.45 0.077 0.468 0.243 ;
        RECT 0.418 0.077 0.468 0.095 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.121 0.18 0.581 0.198 ;
      LAYER M1 ;
        RECT 0.526 0.189 0.576 0.207 ;
        RECT 0.558 0.121 0.576 0.207 ;
        RECT 0.107 0.189 0.144 0.207 ;
        RECT 0.126 0.121 0.144 0.207 ;
      LAYER V1 ;
        RECT 0.126 0.18 0.144 0.198 ;
        RECT 0.558 0.18 0.576 0.198 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 0.092 0.225 0.193 0.243 ;
      RECT 0.174 0.189 0.193 0.243 ;
      RECT 0.174 0.189 0.414 0.207 ;
      RECT 0.396 0.121 0.414 0.207 ;
      RECT 0.174 0.082 0.192 0.243 ;
      RECT 0.256 0.027 0.608 0.045 ;
  END
END XNOR2x1_ASAP7_75t_L

MACRO XNOR2x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x2_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.225 0.44 0.243 ;
        RECT 0.422 0.126 0.44 0.243 ;
        RECT 0.391 0.126 0.44 0.144 ;
        RECT 0.261 0.183 0.279 0.243 ;
        RECT 0.126 0.183 0.279 0.201 ;
        RECT 0.126 0.12 0.144 0.201 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.189 0.38 0.207 ;
        RECT 0.342 0.107 0.36 0.207 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.225 0.576 0.243 ;
        RECT 0.558 0.027 0.576 0.243 ;
        RECT 0.472 0.027 0.576 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.225 0.063 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.477 0.063 0.495 0.151 ;
      RECT 0.423 0.063 0.495 0.081 ;
      RECT 0.423 0.027 0.441 0.081 ;
      RECT 0.018 0.027 0.441 0.045 ;
      RECT 0.302 0.063 0.32 0.195 ;
      RECT 0.072 0.063 0.09 0.149 ;
      RECT 0.072 0.063 0.392 0.081 ;
      RECT 0.099 0.225 0.23 0.243 ;
  END
END XNOR2x2_ASAP7_75t_L

MACRO XNOR2xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.063 0.36 0.164 ;
        RECT 0.207 0.063 0.36 0.081 ;
        RECT 0.207 0.027 0.225 0.081 ;
        RECT 0.072 0.027 0.225 0.045 ;
        RECT 0.072 0.027 0.09 0.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.07 0.144 0.2 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.423 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.225 0.18 0.243 ;
      RECT 0.162 0.075 0.18 0.243 ;
      RECT 0.162 0.189 0.414 0.207 ;
      RECT 0.396 0.121 0.414 0.207 ;
      RECT 0.261 0.027 0.387 0.045 ;
  END
END XNOR2xp5_ASAP7_75t_L

MACRO XOR2x1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x1_ASAP7_75t_L 0 0 ;
  SIZE 0.648 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.298 0.18 0.527 0.198 ;
      LAYER M1 ;
        RECT 0.504 0.118 0.522 0.2 ;
        RECT 0.305 0.126 0.365 0.144 ;
        RECT 0.213 0.185 0.323 0.203 ;
        RECT 0.305 0.126 0.323 0.203 ;
        RECT 0.018 0.225 0.231 0.243 ;
        RECT 0.213 0.185 0.231 0.243 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.034 0.036 0.243 ;
      LAYER V1 ;
        RECT 0.305 0.18 0.323 0.198 ;
        RECT 0.504 0.18 0.522 0.198 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.648 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.027 0.612 0.045 ;
        RECT 0.418 0.175 0.468 0.193 ;
        RECT 0.45 0.027 0.468 0.193 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.121 0.072 0.581 0.09 ;
      LAYER M1 ;
        RECT 0.558 0.063 0.576 0.149 ;
        RECT 0.526 0.063 0.576 0.081 ;
        RECT 0.126 0.063 0.144 0.149 ;
        RECT 0.107 0.063 0.144 0.081 ;
      LAYER V1 ;
        RECT 0.126 0.072 0.144 0.09 ;
        RECT 0.558 0.072 0.576 0.09 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.174 0.027 0.192 0.188 ;
      RECT 0.396 0.063 0.414 0.149 ;
      RECT 0.174 0.063 0.414 0.081 ;
      RECT 0.174 0.027 0.193 0.081 ;
      RECT 0.092 0.027 0.193 0.045 ;
      RECT 0.256 0.225 0.608 0.243 ;
  END
END XOR2x1_ASAP7_75t_L

MACRO XOR2x2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x2_ASAP7_75t_L 0 0 ;
  SIZE 0.594 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.063 0.38 0.081 ;
        RECT 0.342 0.063 0.36 0.163 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.422 0.027 0.44 0.163 ;
        RECT 0.391 0.126 0.44 0.144 ;
        RECT 0.261 0.027 0.44 0.045 ;
        RECT 0.126 0.069 0.279 0.087 ;
        RECT 0.261 0.027 0.279 0.087 ;
        RECT 0.126 0.069 0.144 0.15 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.594 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.225 0.576 0.243 ;
        RECT 0.558 0.027 0.576 0.243 ;
        RECT 0.472 0.027 0.576 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.018 0.225 0.441 0.243 ;
      RECT 0.423 0.189 0.441 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.423 0.189 0.495 0.207 ;
      RECT 0.477 0.119 0.495 0.207 ;
      RECT 0.018 0.027 0.063 0.045 ;
      RECT 0.072 0.189 0.392 0.207 ;
      RECT 0.302 0.075 0.32 0.207 ;
      RECT 0.072 0.121 0.09 0.207 ;
      RECT 0.099 0.027 0.23 0.045 ;
  END
END XOR2x2_ASAP7_75t_L

MACRO XOR2xp5_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2xp5_ASAP7_75t_L 0 0 ;
  SIZE 0.486 BY 0.27 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.189 0.36 0.207 ;
        RECT 0.342 0.12 0.36 0.207 ;
        RECT 0.018 0.225 0.225 0.243 ;
        RECT 0.207 0.189 0.225 0.243 ;
        RECT 0.018 0.126 0.078 0.144 ;
        RECT 0.018 0.034 0.036 0.243 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.106 0.189 0.144 0.207 ;
        RECT 0.126 0.063 0.144 0.207 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 0.486 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.225 0.468 0.243 ;
        RECT 0.45 0.027 0.468 0.243 ;
        RECT 0.256 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.162 0.027 0.18 0.195 ;
      RECT 0.396 0.063 0.414 0.149 ;
      RECT 0.162 0.063 0.414 0.081 ;
      RECT 0.094 0.027 0.18 0.045 ;
      RECT 0.256 0.225 0.387 0.243 ;
  END
END XOR2xp5_ASAP7_75t_L

END LIBRARY
