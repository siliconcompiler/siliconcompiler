VERSION 5.4 ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

MANUFACTURINGGRID 0.01000 ;

MACRO RAM
    CLASS INOUT ;
    FOREIGN RAM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.000 BY 50.000 ;
    SYMMETRY R90 ;
END RAM

END LIBRARY