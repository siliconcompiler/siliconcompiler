module interposer (
    inout [53:0] ios0
);

endmodule
