VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_32x2048_1rw
  FOREIGN sram_32x2048_1rw 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 190.760 BY 313.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.965 0.070 49.035 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.365 0.070 57.435 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.865 0.070 88.935 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.665 0.070 91.735 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.265 0.070 97.335 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.065 0.070 100.135 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.865 0.070 102.935 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.665 0.070 105.735 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.465 0.070 108.535 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.265 0.070 111.335 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.065 0.070 114.135 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.865 0.070 116.935 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.665 0.070 119.735 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.465 0.070 122.535 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.265 0.070 125.335 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.065 0.070 128.135 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.865 0.070 130.935 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.665 0.070 133.735 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.465 0.070 136.535 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.265 0.070 139.335 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.065 0.070 142.135 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.865 0.070 144.935 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.665 0.070 147.735 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.465 0.070 150.535 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.265 0.070 153.335 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.065 0.070 156.135 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.865 0.070 158.935 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.665 0.070 161.735 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.465 0.070 164.535 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.265 0.070 167.335 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.065 0.070 170.135 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.865 0.070 172.935 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.665 0.070 175.735 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.365 0.070 176.435 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.165 0.070 179.235 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.965 0.070 182.035 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.765 0.070 184.835 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.565 0.070 187.635 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.365 0.070 190.435 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.165 0.070 193.235 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.965 0.070 196.035 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.765 0.070 198.835 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.565 0.070 201.635 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.365 0.070 204.435 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.165 0.070 207.235 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.965 0.070 210.035 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.765 0.070 212.835 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.565 0.070 215.635 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.365 0.070 218.435 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.165 0.070 221.235 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.965 0.070 224.035 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.765 0.070 226.835 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.565 0.070 229.635 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.365 0.070 232.435 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.165 0.070 235.235 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.965 0.070 238.035 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.765 0.070 240.835 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.565 0.070 243.635 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.365 0.070 246.435 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.165 0.070 249.235 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.965 0.070 252.035 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.765 0.070 254.835 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.565 0.070 257.635 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.365 0.070 260.435 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.165 0.070 263.235 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.865 0.070 263.935 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.665 0.070 266.735 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.465 0.070 269.535 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.265 0.070 272.335 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.065 0.070 275.135 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.865 0.070 277.935 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.665 0.070 280.735 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.465 0.070 283.535 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.265 0.070 286.335 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.065 0.070 289.135 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.865 0.070 291.935 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.565 0.070 292.635 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.365 0.070 295.435 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.165 0.070 298.235 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 312.200 ;
      RECT 3.500 1.400 3.780 312.200 ;
      RECT 5.740 1.400 6.020 312.200 ;
      RECT 7.980 1.400 8.260 312.200 ;
      RECT 10.220 1.400 10.500 312.200 ;
      RECT 12.460 1.400 12.740 312.200 ;
      RECT 14.700 1.400 14.980 312.200 ;
      RECT 16.940 1.400 17.220 312.200 ;
      RECT 19.180 1.400 19.460 312.200 ;
      RECT 21.420 1.400 21.700 312.200 ;
      RECT 23.660 1.400 23.940 312.200 ;
      RECT 25.900 1.400 26.180 312.200 ;
      RECT 28.140 1.400 28.420 312.200 ;
      RECT 30.380 1.400 30.660 312.200 ;
      RECT 32.620 1.400 32.900 312.200 ;
      RECT 34.860 1.400 35.140 312.200 ;
      RECT 37.100 1.400 37.380 312.200 ;
      RECT 39.340 1.400 39.620 312.200 ;
      RECT 41.580 1.400 41.860 312.200 ;
      RECT 43.820 1.400 44.100 312.200 ;
      RECT 46.060 1.400 46.340 312.200 ;
      RECT 48.300 1.400 48.580 312.200 ;
      RECT 50.540 1.400 50.820 312.200 ;
      RECT 52.780 1.400 53.060 312.200 ;
      RECT 55.020 1.400 55.300 312.200 ;
      RECT 57.260 1.400 57.540 312.200 ;
      RECT 59.500 1.400 59.780 312.200 ;
      RECT 61.740 1.400 62.020 312.200 ;
      RECT 63.980 1.400 64.260 312.200 ;
      RECT 66.220 1.400 66.500 312.200 ;
      RECT 68.460 1.400 68.740 312.200 ;
      RECT 70.700 1.400 70.980 312.200 ;
      RECT 72.940 1.400 73.220 312.200 ;
      RECT 75.180 1.400 75.460 312.200 ;
      RECT 77.420 1.400 77.700 312.200 ;
      RECT 79.660 1.400 79.940 312.200 ;
      RECT 81.900 1.400 82.180 312.200 ;
      RECT 84.140 1.400 84.420 312.200 ;
      RECT 86.380 1.400 86.660 312.200 ;
      RECT 88.620 1.400 88.900 312.200 ;
      RECT 90.860 1.400 91.140 312.200 ;
      RECT 93.100 1.400 93.380 312.200 ;
      RECT 95.340 1.400 95.620 312.200 ;
      RECT 97.580 1.400 97.860 312.200 ;
      RECT 99.820 1.400 100.100 312.200 ;
      RECT 102.060 1.400 102.340 312.200 ;
      RECT 104.300 1.400 104.580 312.200 ;
      RECT 106.540 1.400 106.820 312.200 ;
      RECT 108.780 1.400 109.060 312.200 ;
      RECT 111.020 1.400 111.300 312.200 ;
      RECT 113.260 1.400 113.540 312.200 ;
      RECT 115.500 1.400 115.780 312.200 ;
      RECT 117.740 1.400 118.020 312.200 ;
      RECT 119.980 1.400 120.260 312.200 ;
      RECT 122.220 1.400 122.500 312.200 ;
      RECT 124.460 1.400 124.740 312.200 ;
      RECT 126.700 1.400 126.980 312.200 ;
      RECT 128.940 1.400 129.220 312.200 ;
      RECT 131.180 1.400 131.460 312.200 ;
      RECT 133.420 1.400 133.700 312.200 ;
      RECT 135.660 1.400 135.940 312.200 ;
      RECT 137.900 1.400 138.180 312.200 ;
      RECT 140.140 1.400 140.420 312.200 ;
      RECT 142.380 1.400 142.660 312.200 ;
      RECT 144.620 1.400 144.900 312.200 ;
      RECT 146.860 1.400 147.140 312.200 ;
      RECT 149.100 1.400 149.380 312.200 ;
      RECT 151.340 1.400 151.620 312.200 ;
      RECT 153.580 1.400 153.860 312.200 ;
      RECT 155.820 1.400 156.100 312.200 ;
      RECT 158.060 1.400 158.340 312.200 ;
      RECT 160.300 1.400 160.580 312.200 ;
      RECT 162.540 1.400 162.820 312.200 ;
      RECT 164.780 1.400 165.060 312.200 ;
      RECT 167.020 1.400 167.300 312.200 ;
      RECT 169.260 1.400 169.540 312.200 ;
      RECT 171.500 1.400 171.780 312.200 ;
      RECT 173.740 1.400 174.020 312.200 ;
      RECT 175.980 1.400 176.260 312.200 ;
      RECT 178.220 1.400 178.500 312.200 ;
      RECT 180.460 1.400 180.740 312.200 ;
      RECT 182.700 1.400 182.980 312.200 ;
      RECT 184.940 1.400 185.220 312.200 ;
      RECT 187.180 1.400 187.460 312.200 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 312.200 ;
      RECT 4.620 1.400 4.900 312.200 ;
      RECT 6.860 1.400 7.140 312.200 ;
      RECT 9.100 1.400 9.380 312.200 ;
      RECT 11.340 1.400 11.620 312.200 ;
      RECT 13.580 1.400 13.860 312.200 ;
      RECT 15.820 1.400 16.100 312.200 ;
      RECT 18.060 1.400 18.340 312.200 ;
      RECT 20.300 1.400 20.580 312.200 ;
      RECT 22.540 1.400 22.820 312.200 ;
      RECT 24.780 1.400 25.060 312.200 ;
      RECT 27.020 1.400 27.300 312.200 ;
      RECT 29.260 1.400 29.540 312.200 ;
      RECT 31.500 1.400 31.780 312.200 ;
      RECT 33.740 1.400 34.020 312.200 ;
      RECT 35.980 1.400 36.260 312.200 ;
      RECT 38.220 1.400 38.500 312.200 ;
      RECT 40.460 1.400 40.740 312.200 ;
      RECT 42.700 1.400 42.980 312.200 ;
      RECT 44.940 1.400 45.220 312.200 ;
      RECT 47.180 1.400 47.460 312.200 ;
      RECT 49.420 1.400 49.700 312.200 ;
      RECT 51.660 1.400 51.940 312.200 ;
      RECT 53.900 1.400 54.180 312.200 ;
      RECT 56.140 1.400 56.420 312.200 ;
      RECT 58.380 1.400 58.660 312.200 ;
      RECT 60.620 1.400 60.900 312.200 ;
      RECT 62.860 1.400 63.140 312.200 ;
      RECT 65.100 1.400 65.380 312.200 ;
      RECT 67.340 1.400 67.620 312.200 ;
      RECT 69.580 1.400 69.860 312.200 ;
      RECT 71.820 1.400 72.100 312.200 ;
      RECT 74.060 1.400 74.340 312.200 ;
      RECT 76.300 1.400 76.580 312.200 ;
      RECT 78.540 1.400 78.820 312.200 ;
      RECT 80.780 1.400 81.060 312.200 ;
      RECT 83.020 1.400 83.300 312.200 ;
      RECT 85.260 1.400 85.540 312.200 ;
      RECT 87.500 1.400 87.780 312.200 ;
      RECT 89.740 1.400 90.020 312.200 ;
      RECT 91.980 1.400 92.260 312.200 ;
      RECT 94.220 1.400 94.500 312.200 ;
      RECT 96.460 1.400 96.740 312.200 ;
      RECT 98.700 1.400 98.980 312.200 ;
      RECT 100.940 1.400 101.220 312.200 ;
      RECT 103.180 1.400 103.460 312.200 ;
      RECT 105.420 1.400 105.700 312.200 ;
      RECT 107.660 1.400 107.940 312.200 ;
      RECT 109.900 1.400 110.180 312.200 ;
      RECT 112.140 1.400 112.420 312.200 ;
      RECT 114.380 1.400 114.660 312.200 ;
      RECT 116.620 1.400 116.900 312.200 ;
      RECT 118.860 1.400 119.140 312.200 ;
      RECT 121.100 1.400 121.380 312.200 ;
      RECT 123.340 1.400 123.620 312.200 ;
      RECT 125.580 1.400 125.860 312.200 ;
      RECT 127.820 1.400 128.100 312.200 ;
      RECT 130.060 1.400 130.340 312.200 ;
      RECT 132.300 1.400 132.580 312.200 ;
      RECT 134.540 1.400 134.820 312.200 ;
      RECT 136.780 1.400 137.060 312.200 ;
      RECT 139.020 1.400 139.300 312.200 ;
      RECT 141.260 1.400 141.540 312.200 ;
      RECT 143.500 1.400 143.780 312.200 ;
      RECT 145.740 1.400 146.020 312.200 ;
      RECT 147.980 1.400 148.260 312.200 ;
      RECT 150.220 1.400 150.500 312.200 ;
      RECT 152.460 1.400 152.740 312.200 ;
      RECT 154.700 1.400 154.980 312.200 ;
      RECT 156.940 1.400 157.220 312.200 ;
      RECT 159.180 1.400 159.460 312.200 ;
      RECT 161.420 1.400 161.700 312.200 ;
      RECT 163.660 1.400 163.940 312.200 ;
      RECT 165.900 1.400 166.180 312.200 ;
      RECT 168.140 1.400 168.420 312.200 ;
      RECT 170.380 1.400 170.660 312.200 ;
      RECT 172.620 1.400 172.900 312.200 ;
      RECT 174.860 1.400 175.140 312.200 ;
      RECT 177.100 1.400 177.380 312.200 ;
      RECT 179.340 1.400 179.620 312.200 ;
      RECT 181.580 1.400 181.860 312.200 ;
      RECT 183.820 1.400 184.100 312.200 ;
      RECT 186.060 1.400 186.340 312.200 ;
      RECT 188.300 1.400 188.580 312.200 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 190.760 313.600 ;
    LAYER metal2 ;
    RECT 0 0 190.760 313.600 ;
    LAYER metal3 ;
    RECT 0.070 0 190.760 313.600 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 4.165 ;
    RECT 0 4.235 0.070 6.965 ;
    RECT 0 7.035 0.070 9.765 ;
    RECT 0 9.835 0.070 12.565 ;
    RECT 0 12.635 0.070 15.365 ;
    RECT 0 15.435 0.070 18.165 ;
    RECT 0 18.235 0.070 20.965 ;
    RECT 0 21.035 0.070 23.765 ;
    RECT 0 23.835 0.070 26.565 ;
    RECT 0 26.635 0.070 29.365 ;
    RECT 0 29.435 0.070 32.165 ;
    RECT 0 32.235 0.070 34.965 ;
    RECT 0 35.035 0.070 37.765 ;
    RECT 0 37.835 0.070 40.565 ;
    RECT 0 40.635 0.070 43.365 ;
    RECT 0 43.435 0.070 46.165 ;
    RECT 0 46.235 0.070 48.965 ;
    RECT 0 49.035 0.070 51.765 ;
    RECT 0 51.835 0.070 54.565 ;
    RECT 0 54.635 0.070 57.365 ;
    RECT 0 57.435 0.070 60.165 ;
    RECT 0 60.235 0.070 62.965 ;
    RECT 0 63.035 0.070 65.765 ;
    RECT 0 65.835 0.070 68.565 ;
    RECT 0 68.635 0.070 71.365 ;
    RECT 0 71.435 0.070 74.165 ;
    RECT 0 74.235 0.070 76.965 ;
    RECT 0 77.035 0.070 79.765 ;
    RECT 0 79.835 0.070 82.565 ;
    RECT 0 82.635 0.070 85.365 ;
    RECT 0 85.435 0.070 88.165 ;
    RECT 0 88.235 0.070 88.865 ;
    RECT 0 88.935 0.070 91.665 ;
    RECT 0 91.735 0.070 94.465 ;
    RECT 0 94.535 0.070 97.265 ;
    RECT 0 97.335 0.070 100.065 ;
    RECT 0 100.135 0.070 102.865 ;
    RECT 0 102.935 0.070 105.665 ;
    RECT 0 105.735 0.070 108.465 ;
    RECT 0 108.535 0.070 111.265 ;
    RECT 0 111.335 0.070 114.065 ;
    RECT 0 114.135 0.070 116.865 ;
    RECT 0 116.935 0.070 119.665 ;
    RECT 0 119.735 0.070 122.465 ;
    RECT 0 122.535 0.070 125.265 ;
    RECT 0 125.335 0.070 128.065 ;
    RECT 0 128.135 0.070 130.865 ;
    RECT 0 130.935 0.070 133.665 ;
    RECT 0 133.735 0.070 136.465 ;
    RECT 0 136.535 0.070 139.265 ;
    RECT 0 139.335 0.070 142.065 ;
    RECT 0 142.135 0.070 144.865 ;
    RECT 0 144.935 0.070 147.665 ;
    RECT 0 147.735 0.070 150.465 ;
    RECT 0 150.535 0.070 153.265 ;
    RECT 0 153.335 0.070 156.065 ;
    RECT 0 156.135 0.070 158.865 ;
    RECT 0 158.935 0.070 161.665 ;
    RECT 0 161.735 0.070 164.465 ;
    RECT 0 164.535 0.070 167.265 ;
    RECT 0 167.335 0.070 170.065 ;
    RECT 0 170.135 0.070 172.865 ;
    RECT 0 172.935 0.070 175.665 ;
    RECT 0 175.735 0.070 176.365 ;
    RECT 0 176.435 0.070 179.165 ;
    RECT 0 179.235 0.070 181.965 ;
    RECT 0 182.035 0.070 184.765 ;
    RECT 0 184.835 0.070 187.565 ;
    RECT 0 187.635 0.070 190.365 ;
    RECT 0 190.435 0.070 193.165 ;
    RECT 0 193.235 0.070 195.965 ;
    RECT 0 196.035 0.070 198.765 ;
    RECT 0 198.835 0.070 201.565 ;
    RECT 0 201.635 0.070 204.365 ;
    RECT 0 204.435 0.070 207.165 ;
    RECT 0 207.235 0.070 209.965 ;
    RECT 0 210.035 0.070 212.765 ;
    RECT 0 212.835 0.070 215.565 ;
    RECT 0 215.635 0.070 218.365 ;
    RECT 0 218.435 0.070 221.165 ;
    RECT 0 221.235 0.070 223.965 ;
    RECT 0 224.035 0.070 226.765 ;
    RECT 0 226.835 0.070 229.565 ;
    RECT 0 229.635 0.070 232.365 ;
    RECT 0 232.435 0.070 235.165 ;
    RECT 0 235.235 0.070 237.965 ;
    RECT 0 238.035 0.070 240.765 ;
    RECT 0 240.835 0.070 243.565 ;
    RECT 0 243.635 0.070 246.365 ;
    RECT 0 246.435 0.070 249.165 ;
    RECT 0 249.235 0.070 251.965 ;
    RECT 0 252.035 0.070 254.765 ;
    RECT 0 254.835 0.070 257.565 ;
    RECT 0 257.635 0.070 260.365 ;
    RECT 0 260.435 0.070 263.165 ;
    RECT 0 263.235 0.070 263.865 ;
    RECT 0 263.935 0.070 266.665 ;
    RECT 0 266.735 0.070 269.465 ;
    RECT 0 269.535 0.070 272.265 ;
    RECT 0 272.335 0.070 275.065 ;
    RECT 0 275.135 0.070 277.865 ;
    RECT 0 277.935 0.070 280.665 ;
    RECT 0 280.735 0.070 283.465 ;
    RECT 0 283.535 0.070 286.265 ;
    RECT 0 286.335 0.070 289.065 ;
    RECT 0 289.135 0.070 291.865 ;
    RECT 0 291.935 0.070 292.565 ;
    RECT 0 292.635 0.070 295.365 ;
    RECT 0 295.435 0.070 298.165 ;
    RECT 0 298.235 0.070 313.600 ;
    LAYER metal4 ;
    RECT 0 0 190.760 1.400 ;
    RECT 0 312.200 190.760 313.600 ;
    RECT 0.000 1.400 1.260 312.200 ;
    RECT 1.540 1.400 2.380 312.200 ;
    RECT 2.660 1.400 3.500 312.200 ;
    RECT 3.780 1.400 4.620 312.200 ;
    RECT 4.900 1.400 5.740 312.200 ;
    RECT 6.020 1.400 6.860 312.200 ;
    RECT 7.140 1.400 7.980 312.200 ;
    RECT 8.260 1.400 9.100 312.200 ;
    RECT 9.380 1.400 10.220 312.200 ;
    RECT 10.500 1.400 11.340 312.200 ;
    RECT 11.620 1.400 12.460 312.200 ;
    RECT 12.740 1.400 13.580 312.200 ;
    RECT 13.860 1.400 14.700 312.200 ;
    RECT 14.980 1.400 15.820 312.200 ;
    RECT 16.100 1.400 16.940 312.200 ;
    RECT 17.220 1.400 18.060 312.200 ;
    RECT 18.340 1.400 19.180 312.200 ;
    RECT 19.460 1.400 20.300 312.200 ;
    RECT 20.580 1.400 21.420 312.200 ;
    RECT 21.700 1.400 22.540 312.200 ;
    RECT 22.820 1.400 23.660 312.200 ;
    RECT 23.940 1.400 24.780 312.200 ;
    RECT 25.060 1.400 25.900 312.200 ;
    RECT 26.180 1.400 27.020 312.200 ;
    RECT 27.300 1.400 28.140 312.200 ;
    RECT 28.420 1.400 29.260 312.200 ;
    RECT 29.540 1.400 30.380 312.200 ;
    RECT 30.660 1.400 31.500 312.200 ;
    RECT 31.780 1.400 32.620 312.200 ;
    RECT 32.900 1.400 33.740 312.200 ;
    RECT 34.020 1.400 34.860 312.200 ;
    RECT 35.140 1.400 35.980 312.200 ;
    RECT 36.260 1.400 37.100 312.200 ;
    RECT 37.380 1.400 38.220 312.200 ;
    RECT 38.500 1.400 39.340 312.200 ;
    RECT 39.620 1.400 40.460 312.200 ;
    RECT 40.740 1.400 41.580 312.200 ;
    RECT 41.860 1.400 42.700 312.200 ;
    RECT 42.980 1.400 43.820 312.200 ;
    RECT 44.100 1.400 44.940 312.200 ;
    RECT 45.220 1.400 46.060 312.200 ;
    RECT 46.340 1.400 47.180 312.200 ;
    RECT 47.460 1.400 48.300 312.200 ;
    RECT 48.580 1.400 49.420 312.200 ;
    RECT 49.700 1.400 50.540 312.200 ;
    RECT 50.820 1.400 51.660 312.200 ;
    RECT 51.940 1.400 52.780 312.200 ;
    RECT 53.060 1.400 53.900 312.200 ;
    RECT 54.180 1.400 55.020 312.200 ;
    RECT 55.300 1.400 56.140 312.200 ;
    RECT 56.420 1.400 57.260 312.200 ;
    RECT 57.540 1.400 58.380 312.200 ;
    RECT 58.660 1.400 59.500 312.200 ;
    RECT 59.780 1.400 60.620 312.200 ;
    RECT 60.900 1.400 61.740 312.200 ;
    RECT 62.020 1.400 62.860 312.200 ;
    RECT 63.140 1.400 63.980 312.200 ;
    RECT 64.260 1.400 65.100 312.200 ;
    RECT 65.380 1.400 66.220 312.200 ;
    RECT 66.500 1.400 67.340 312.200 ;
    RECT 67.620 1.400 68.460 312.200 ;
    RECT 68.740 1.400 69.580 312.200 ;
    RECT 69.860 1.400 70.700 312.200 ;
    RECT 70.980 1.400 71.820 312.200 ;
    RECT 72.100 1.400 72.940 312.200 ;
    RECT 73.220 1.400 74.060 312.200 ;
    RECT 74.340 1.400 75.180 312.200 ;
    RECT 75.460 1.400 76.300 312.200 ;
    RECT 76.580 1.400 77.420 312.200 ;
    RECT 77.700 1.400 78.540 312.200 ;
    RECT 78.820 1.400 79.660 312.200 ;
    RECT 79.940 1.400 80.780 312.200 ;
    RECT 81.060 1.400 81.900 312.200 ;
    RECT 82.180 1.400 83.020 312.200 ;
    RECT 83.300 1.400 84.140 312.200 ;
    RECT 84.420 1.400 85.260 312.200 ;
    RECT 85.540 1.400 86.380 312.200 ;
    RECT 86.660 1.400 87.500 312.200 ;
    RECT 87.780 1.400 88.620 312.200 ;
    RECT 88.900 1.400 89.740 312.200 ;
    RECT 90.020 1.400 90.860 312.200 ;
    RECT 91.140 1.400 91.980 312.200 ;
    RECT 92.260 1.400 93.100 312.200 ;
    RECT 93.380 1.400 94.220 312.200 ;
    RECT 94.500 1.400 95.340 312.200 ;
    RECT 95.620 1.400 96.460 312.200 ;
    RECT 96.740 1.400 97.580 312.200 ;
    RECT 97.860 1.400 98.700 312.200 ;
    RECT 98.980 1.400 99.820 312.200 ;
    RECT 100.100 1.400 100.940 312.200 ;
    RECT 101.220 1.400 102.060 312.200 ;
    RECT 102.340 1.400 103.180 312.200 ;
    RECT 103.460 1.400 104.300 312.200 ;
    RECT 104.580 1.400 105.420 312.200 ;
    RECT 105.700 1.400 106.540 312.200 ;
    RECT 106.820 1.400 107.660 312.200 ;
    RECT 107.940 1.400 108.780 312.200 ;
    RECT 109.060 1.400 109.900 312.200 ;
    RECT 110.180 1.400 111.020 312.200 ;
    RECT 111.300 1.400 112.140 312.200 ;
    RECT 112.420 1.400 113.260 312.200 ;
    RECT 113.540 1.400 114.380 312.200 ;
    RECT 114.660 1.400 115.500 312.200 ;
    RECT 115.780 1.400 116.620 312.200 ;
    RECT 116.900 1.400 117.740 312.200 ;
    RECT 118.020 1.400 118.860 312.200 ;
    RECT 119.140 1.400 119.980 312.200 ;
    RECT 120.260 1.400 121.100 312.200 ;
    RECT 121.380 1.400 122.220 312.200 ;
    RECT 122.500 1.400 123.340 312.200 ;
    RECT 123.620 1.400 124.460 312.200 ;
    RECT 124.740 1.400 125.580 312.200 ;
    RECT 125.860 1.400 126.700 312.200 ;
    RECT 126.980 1.400 127.820 312.200 ;
    RECT 128.100 1.400 128.940 312.200 ;
    RECT 129.220 1.400 130.060 312.200 ;
    RECT 130.340 1.400 131.180 312.200 ;
    RECT 131.460 1.400 132.300 312.200 ;
    RECT 132.580 1.400 133.420 312.200 ;
    RECT 133.700 1.400 134.540 312.200 ;
    RECT 134.820 1.400 135.660 312.200 ;
    RECT 135.940 1.400 136.780 312.200 ;
    RECT 137.060 1.400 137.900 312.200 ;
    RECT 138.180 1.400 139.020 312.200 ;
    RECT 139.300 1.400 140.140 312.200 ;
    RECT 140.420 1.400 141.260 312.200 ;
    RECT 141.540 1.400 142.380 312.200 ;
    RECT 142.660 1.400 143.500 312.200 ;
    RECT 143.780 1.400 144.620 312.200 ;
    RECT 144.900 1.400 145.740 312.200 ;
    RECT 146.020 1.400 146.860 312.200 ;
    RECT 147.140 1.400 147.980 312.200 ;
    RECT 148.260 1.400 149.100 312.200 ;
    RECT 149.380 1.400 150.220 312.200 ;
    RECT 150.500 1.400 151.340 312.200 ;
    RECT 151.620 1.400 152.460 312.200 ;
    RECT 152.740 1.400 153.580 312.200 ;
    RECT 153.860 1.400 154.700 312.200 ;
    RECT 154.980 1.400 155.820 312.200 ;
    RECT 156.100 1.400 156.940 312.200 ;
    RECT 157.220 1.400 158.060 312.200 ;
    RECT 158.340 1.400 159.180 312.200 ;
    RECT 159.460 1.400 160.300 312.200 ;
    RECT 160.580 1.400 161.420 312.200 ;
    RECT 161.700 1.400 162.540 312.200 ;
    RECT 162.820 1.400 163.660 312.200 ;
    RECT 163.940 1.400 164.780 312.200 ;
    RECT 165.060 1.400 165.900 312.200 ;
    RECT 166.180 1.400 167.020 312.200 ;
    RECT 167.300 1.400 168.140 312.200 ;
    RECT 168.420 1.400 169.260 312.200 ;
    RECT 169.540 1.400 170.380 312.200 ;
    RECT 170.660 1.400 171.500 312.200 ;
    RECT 171.780 1.400 172.620 312.200 ;
    RECT 172.900 1.400 173.740 312.200 ;
    RECT 174.020 1.400 174.860 312.200 ;
    RECT 175.140 1.400 175.980 312.200 ;
    RECT 176.260 1.400 177.100 312.200 ;
    RECT 177.380 1.400 178.220 312.200 ;
    RECT 178.500 1.400 179.340 312.200 ;
    RECT 179.620 1.400 180.460 312.200 ;
    RECT 180.740 1.400 181.580 312.200 ;
    RECT 181.860 1.400 182.700 312.200 ;
    RECT 182.980 1.400 183.820 312.200 ;
    RECT 184.100 1.400 184.940 312.200 ;
    RECT 185.220 1.400 186.060 312.200 ;
    RECT 186.340 1.400 187.180 312.200 ;
    RECT 187.460 1.400 188.300 312.200 ;
    RECT 188.580 1.400 190.760 312.200 ;
    LAYER OVERLAP ;
    RECT 0 0 190.760 313.600 ;
  END
END sram_32x2048_1rw

END LIBRARY
