# BSD 3-Clause License
# 
# Copyright 2020 Lawrence T. Clark, Vinay Vashishtha, or Arizona State
# University
# 
# Redistribution and use in source and binary forms, with or without
# modification, are permitted provided that the following conditions are met:
# 
# 1. Redistributions of source code must retain the above copyright notice,
# this list of conditions and the following disclaimer.
# 
# 2. Redistributions in binary form must reproduce the above copyright
# notice, this list of conditions and the following disclaimer in the
# documentation and/or other materials provided with the distribution.
# 
# 3. Neither the name of the copyright holder nor the names of its
# contributors may be used to endorse or promote products derived from this
# software without specific prior written permission.
# 
# THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
# AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
# IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
# ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
# LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
# CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
# SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
# INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
# CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
# ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
# POSSIBILITY OF SUCH DAMAGE.

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS
MANUFACTURINGGRID 0.004 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_PITCH STRING ;
  LAYER LEF58_GAP STRING ;
  LAYER LEF58_EOLKEEPOUT STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_CORNERSPACING STRING ;
  LAYER LEF58_WIDTHTABLE STRING ;
  LAYER LEF58_CUTCLASS STRING ;
  LAYER LEF58_SPACINGTABLE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_RIGHTWAYONGRIDONLY STRING ;
  LAYER LEF58_RECTONLY STRING ;
END PROPERTYDEFINITIONS

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER Gate
  TYPE MASTERSLICE ;
END Gate

LAYER Active
  TYPE MASTERSLICE ;
END Active

LAYER V0
  TYPE CUT ;
  SPACING 0.072 ;
  WIDTH 0.072 ;
END V0

LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.144 ;
  WIDTH 0.072 ;
  SPACING 0.072 ;
  AREA 0.010656 ;                   # Min Area # This should ideally be 16x not 4x as each dimension is scaled up by 16
                                    # we only allow landing on pins (set in router) so area should not matter
  SPACING 0.072 RANGE 0.144 4.000 ; # This rule is redundant with the SPACING rule

  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.073 EXTENSION 0 0 0.124 ;" ; #  Tip to Tip Spacing

  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERONLY 0.040 WIDTH 0.072 SPACING 0.072 ;" ; 
OFFSET 0.0 ;

END M1

LAYER V1
  TYPE CUT ;
  SPACING 0.072 ;     # unlike generate, this is really spacing, not center to center.
  WIDTH 0.072 ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.072 ; # Min Width
  SPACING 0.072 ; # Min Spacing

  OFFSET -1.080 ;

  #  MINSIZE is set so that the minimum lenght of a segment is 36nm. At the proper rule size of
  #  31nm, the lines can't be minimum space. This causes DRCs (like crazy). Same for M3
  #  MINSIZE 0.112 0.072 ; 
  # area is adjusted to match this (Nanoroute requires both AREA and MINSIZE)

  AREA 0.010656 ;
  MINSIZE 0.148 0.072 ; 

  PITCH 0.180 0.144 ;

  # this enforces the correct routing tracks on M2 with wide M2 power rails

  PROPERTY LEF58_PITCH "
   PITCH 0.144 FIRSTLASTPITCH 0.180 
   ;
  " ;

  # this checks for distance in any direction so is not correct
  # 0.070 is to avoid conflicts with the adjacent lines. This should be caught by CORNERSPACING below
  #   SPACING 0.124 ENDOFLINE 0.1 WITHIN 0.070 ;

  PROPERTY LEF58_SPACING 
    " SPACING 0.072 ENDOFLINE 0.1 WITHIN 0.08 ENDTOEND 0.124 
      PARALLELEDGE 0.100 WITHIN 0.08 ; " ;	   

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.1 EXTENSION 0.0 0.05 0.124 CORNERONLY ;
  " ;

  PROPERTY LEF58_CORNERSPACING "
     CORNERSPACING CONVEXCORNER WIDTH 0.000 SPACING 0.080 ;
  " ; # CORNER to CORNER SPACING Rule

  # Originally no width table for M2 since it is the follow rails. 
  # They can be 1x or 2x (2x causes DRCs on SAV V1). However, this seems to allow a double width M2
  # on vias, which violates. Thus, this is added. Note that wide power follow rails will violate.

  PROPERTY LEF58_WIDTHTABLE "
      WIDTHTABLE 0.072 0.36 0.648 0.936 1.224 1.512 ; 
  " ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M2

LAYER V2
  TYPE CUT ;
  SPACING 0.072 ;
  WIDTH 0.072 ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.144 ;
  OFFSET 0.0 ;
  WIDTH 0.072 ; # Min Width
  SPACING 0.072 ; # Min Spacing

  #  MINSIZE is set so that the minimum lenght of a segment is 36nm. At the proper rule size of
  #  31nm, the lines can't be minimum space. This causes DRCs (like crazy). Same for M2
  #  MINSIZE 0.112 0.072 ; 
  # area is adjusted to match this (Nanoroute requires both AREA and MINSIZE)

  AREA 0.010656 ;
  MINSIZE 0.148 0.072 ; 

  PROPERTY LEF58_SPACING 
    " SPACING 0.072 ENDOFLINE 0.1 WITHIN 0.05 ENDTOEND 0.124  
      PARALLELEDGE 0.100 WITHIN 0.08 ; " ;	  

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.1 EXTENSION 0.0 0.05 0.124 CORNERONLY ;
  " ;

  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.000 SPACING 0.080 
   ;
  " ; # CORNER to CORNER SPACING Rule

  # to make the special route widths integer values of the tracks, i.e., 1, 5, 9, 13... min widths
  # the widths should be calculated in the APR tool, since viaGen does not seem to respect these

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.072 0.36 0.648 0.936 1.224 1.512 ; " ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M3

LAYER V3
  TYPE CUT ;
#  SPACING 0.072 ;
#  WIDTH 0.072 ;

  # different format to allow long vias for SAV power connections

  PROPERTY LEF58_CUTCLASS "  
    CUTCLASS V3       WIDTH 0.072 LENGTH 0.096 CUTS 1  ; 
    CUTCLASS V3_0p480 WIDTH 0.072 LENGTH 0.480 CUTS 4  ;
    CUTCLASS V3_0p864 WIDTH 0.072 LENGTH 0.864 CUTS 8  ;
  " ;

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      DEFAULT 0.136
      CUTCLASS   V3 V3_0p480 V3_0p864
        V3       -  -        -        -  - -
        V3_0p480 -  -        -        -  - -
        V3_0p864 -  -        -        -  - -
    ;
  " ;

#   ENCLOSURE CUTCLASS V3 END 0.02 SIDE 0.0 ;
  # covered below? 
  # ENCLOSURE CUTCLASS V3       END 0.02 SIDE 0.0 ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS V3 BELOW EOL 0.0 0.020 0.0 ;
    ENCLOSURE CUTCLASS V3 ABOVE EOL 0.0 0.044 0.0 ;
    ENCLOSURE CUTCLASS V3_0p480 END 0.0  SIDE 0.0 ;
    ENCLOSURE CUTCLASS V3_0p864 END 0.0  SIDE 0.0 ;
  " ;

END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.192 ;
  WIDTH 0.096 ;
  SPACING 0.096 ;

  OFFSET 0.012 ;

  AREA 0.032 ; 

  PROPERTY LEF58_SPACING "
    SPACING 0.096 ENDOFLINE 0.1 WITHIN 0.160 ENDTOEND 0.160 ; " ;	  

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.096 0.480 0.864 1.248 1.632 ; " ;

  PROPERTY LEF58_CORNERSPACING "
    CORNERSPACING CONVEXCORNER CORNERONLY 0.192
      WIDTH 0.000 SPACING 0.160 ;
  " ;

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.1 EXTENSION 0.192 0.097 0.192 CORNERONLY ;
  " ;

  # spacing table is required for the rule that has wide metal requires a 72nm (288 scaled)
  # spacing between wide and minimum metals 

  SPACINGTABLE
    PARALLELRUNLENGTH 0.00
      WIDTH 0.000     0.096
      WIDTH 0.100     0.288 ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M4

LAYER V4
  TYPE CUT ;

  # spacing is 4 * 34 = 136
  # SPACING 0.136 ;
  # WIDTH 0.072 ;
  # ENCLOSURE 0.044 0.0 ;

  PROPERTY LEF58_CUTCLASS "  
    CUTCLASS Vx       WIDTH 0.096 LENGTH 0.096 ; 
    CUTCLASS Vx_0p480 WIDTH 0.096 LENGTH 0.480 CUTS 4  ;
    CUTCLASS Vx_0p864 WIDTH 0.096 LENGTH 0.864 CUTS 8  ;
    CUTCLASS Vx_1p248 WIDTH 0.096 LENGTH 1.248 CUTS 12 ;
    CUTCLASS Vx_1p632 WIDTH 0.096 LENGTH 1.632 CUTS 16 ;
  " ;

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      DEFAULT 0.136
      CUTCLASS   Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
        Vx       -  -        -        -        - -  -        -        -        -
        Vx_0p480 -  -        -        -        - -  -        -        -        -
	Vx_0p864 -  -        -        -        - -  -        -        -        -
	Vx_1p248 -  -        -        -        - -  -        -        -        -
	Vx_1p632 -  -        -        -        - -  -        -        -        -
    ;
  " ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS Vx 0.044 0.0 ;
    ENCLOSURE CUTCLASS Vx EOL   0.0 0.044 0.044 ;
    ENCLOSURE CUTCLASS Vx_0p480 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_0p864 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_1p248 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_1p632 END 0.00 SIDE 0.0 ;
  " ;

END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.192 ;
  WIDTH 0.096 ;
  SPACING 0.096 ;
  OFFSET 0.0 ;

  AREA 0.032 ; 

  PROPERTY LEF58_SPACING "
    SPACING 0.096 ENDOFLINE 0.1 WITHIN 0.160 ENDTOEND 0.160 ; " ;	  

  MINIMUMDENSITY 60 ;
  MAXIMUMDENSITY 360 ;
  DENSITYCHECKWINDOW 80 80 ;
  DENSITYCHECKSTEP 40 ;

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.096 0.480 0.864 1.248 1.632 2.016 2.400 2.784 3.168 3.552 3.936 ; " ;

  PROPERTY LEF58_CORNERSPACING "
    CORNERSPACING CONVEXCORNER CORNERONLY 0.192
      WIDTH 0.000 SPACING 0.160 ;
  " ;

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.1 EXTENSION 0.192 0.097 0.192
    CORNERONLY ;
  " ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0.00
      WIDTH 0.000     0.096
      WIDTH 0.100     0.288 ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M5

LAYER V5
  TYPE CUT ;

  PROPERTY LEF58_CUTCLASS "  
    CUTCLASS Vx       WIDTH 0.096 LENGTH 0.128 ; 
    CUTCLASS Vx_0p480 WIDTH 0.096 LENGTH 0.640 CUTS 4  ;
    CUTCLASS Vx_0p864 WIDTH 0.096 LENGTH 1.152 CUTS 8  ;
    CUTCLASS Vx_1p248 WIDTH 0.096 LENGTH 1.664 CUTS 12 ;
    CUTCLASS Vx_1p632 WIDTH 0.096 LENGTH 2.176 CUTS 16 ;
  " ;

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      DEFAULT 0.136
      CUTCLASS   Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
        Vx       -  -        -        -        - -  -        -        -        -
        Vx_0p480 -  -        -        -        - -  -        -        -        -
	Vx_0p864 -  -        -        -        - -  -        -        -        -
	Vx_1p248 -  -        -        -        - -  -        -        -        -
	Vx_1p632 -  -        -        -        - -  -        -        -        -
    ;
  " ;

  # end refers to the end of the VIA! Thus, since it is rectangular the proper
  # enclosure is on the side not the end...
  # ENCLOSURE CUTCLASS Vx END 0.0 SIDE 0.044 ;  But--this refers to top and bottom
  # actually passing the rule is done by having the correct vias below.

  PROPERTY LEF58_ENCLOSURE "
  ENCLOSURE CUTCLASS Vx EOL 0.0 0.044 0.044 ;
  ENCLOSURE CUTCLASS Vx_0p480 END 0.00 SIDE 0.0 ;
  ENCLOSURE CUTCLASS Vx_0p864 END 0.00 SIDE 0.0 ;
  ENCLOSURE CUTCLASS Vx_1p248 END 0.00 SIDE 0.0 ;
  ENCLOSURE CUTCLASS Vx_1p632 END 0.00 SIDE 0.0 ;
  " ;

#  PROPERTY LEF58_ENCLOSURE "
#  ENCLOSURE CUTCLASS Vx EOL 0.0 0.044 0.0 ;
#  " ;

END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.256 ;
  WIDTH 0.128 ;
  SPACING 0.128 ;

  AREA 0.035 ;   # Areas still need tweaking

  PROPERTY LEF58_SPACING 
    " SPACING 0.128 ENDOFLINE 0.15 WITHIN 0.160 ENDTOEND 0.160 ; " ;	   

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.128 0.640 1.152 1.664 2.176 ; " ;

  PROPERTY LEF58_CORNERSPACING "
    CORNERSPACING CONVEXCORNER CORNERONLY 0.192
      WIDTH 0.000 SPACING 0.160 ;
  " ;

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.2 EXTENSION 0.192 0.129 0.192 CORNERONLY ;
  " ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0.00
      WIDTH 0.000     0.096
      WIDTH 0.100     0.288 ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M6

LAYER V6
  TYPE CUT ;

  PROPERTY LEF58_CUTCLASS "  
    CUTCLASS Vx       WIDTH 0.128 LENGTH 0.128 ; 
    CUTCLASS Vx_0p640 WIDTH 0.128 LENGTH 0.640 CUTS 4  ;
    CUTCLASS Vx_1p152 WIDTH 0.128 LENGTH 1.152 CUTS 8  ;
    CUTCLASS Vx_1p664 WIDTH 0.128 LENGTH 1.664 CUTS 12 ;
    CUTCLASS Vx_2p176 WIDTH 0.128 LENGTH 2.176 CUTS 16 ;
  " ;

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      DEFAULT 0.136
      CUTCLASS   Vx Vx_0p640 Vx_1p152 Vx_1p664 Vx_2p176
        Vx       -  -        -        -        - -  -        -        -        -
        Vx_0p640 -  -        -        -        - -  -        -        -        -
	Vx_1p152 -  -        -        -        - -  -        -        -        -
	Vx_1p664 -  -        -        -        - -  -        -        -        -
	Vx_2p176 -  -        -        -        - -  -        -        -        -
    ;
  " ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS Vx 0.044  0.0 ;
    ENCLOSURE CUTCLASS Vx EOL 0.0 0.044 0.044 ;
    ENCLOSURE CUTCLASS Vx_0p640 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_1p152 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_1p664 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_2p176 END 0.00 SIDE 0.0 ;
  " ;

END V6

LAYER M7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.256 ;
  WIDTH 0.128 ;
  SPACING 0.128 ;

  AREA 0.035 ;   # Areas still need tweaking

  PROPERTY LEF58_SPACING 
    " SPACING 0.120 ENDOFLINE 0.15 WITHIN 0.160 ENDTOEND 0.160 ; " ;	   

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.128 0.640 1.152 1.664 2.176 ; " ;
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PROPERTY LEF58_CORNERSPACING "
    CORNERSPACING CONVEXCORNER CORNERONLY 0.300
      WIDTH 0.000 SPACING 0.160 ;
  " ;

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.2 EXTENSION 0.192 0.129 0.192
    CORNERONLY ;
  " ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0.00
      WIDTH 0.000     0.096
      WIDTH 0.100     0.288 ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M7

LAYER V7
  TYPE CUT ;
  SPACING 0.184 ;
  WIDTH 0.128 ;
END V7

LAYER M8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.32 0.32 ;
  WIDTH 0.16 ;
  AREA 30.08 ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0 1.599 4.799 7.199 
    WIDTH 0 0.16 0.16 0.16 0.16 
    WIDTH 0.239 0.16 0.16 0.16 0.16 
    WIDTH 0.319 0.16 0.16 0.16 0.16 
    WIDTH 0.479 0.16 0.16 0.16 0.16 
    WIDTH 1.999 0.16 0.16 0.16 2 
    WIDTH 3.999 0.16 0.16 0.16 4 ;

  MINIMUMCUT 2 WIDTH 7.22 WITHIN 6.82 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 7.22 WITHIN 6.82 FROMABOVE ;
  MAXWIDTH 8 ;
  MINSTEP 0.16 STEP ;
END M8

LAYER V8
  TYPE CUT ;
  SPACING 0.228 ;
  WIDTH 0.16 ;
END V8


LAYER M9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.32 0.32 ;
  WIDTH 0.16 ;
  AREA 30.08 ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0 1.599 4.799 7.199 
    WIDTH 0 0.16 0.16 0.16 0.16 
    WIDTH 0.239 0.16 0.16 0.16 0.16 
    WIDTH 0.319 0.16 0.16 0.16 0.16 
    WIDTH 0.479 0.16 0.16 0.16 0.16 
    WIDTH 1.999 0.16 0.16 0.16 2 
    WIDTH 3.999 0.16 0.16 0.16 4 ;

  MINIMUMCUT 2 WIDTH 7.22 WITHIN 6.82 FROMABOVE ;
  MINSTEP 0.16 STEP ;
END M9

LAYER V9
  TYPE CUT ;
  SPACING 0.228 ;
  WIDTH 0.16 ;
END V9

LAYER Pad
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.32 0.32 ;
  WIDTH 0.16 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 47.999 
    WIDTH 0 8 8 
    WIDTH 47.999 8 12 ;
  MINIMUMCUT 1 WIDTH 0.16 WITHIN 6.82 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 1.44 WITHIN 6.82 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 7.22 WITHIN 6.82 FROMBELOW ;
  MINIMUMDENSITY 80 ;
  MAXIMUMDENSITY 320 ;
  DENSITYCHECKWINDOW 400 400 ;
  DENSITYCHECKSTEP 200 ;
END Pad

# vias

VIA VIA9Pad Default
  LAYER M9 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER Pad ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER V9 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END VIA9Pad

VIA VIA89 Default
  LAYER M8 ;
    RECT -0.08 -0.08 0.08 0.08 ;
  LAYER M9 ;
    RECT -0.08 -0.08 0.08 0.08 ;
  LAYER V8 ;
    RECT -0.08 -0.08 0.08 0.08 ;
END VIA89

VIA VIA78 Default
  LAYER M7 ;
    RECT -0.064 -0.108 0.064 0.108 ;
  LAYER M8 ;
    RECT -0.108 -0.064 0.108 0.064 ;
  LAYER V7 ;
    RECT -0.064 -0.064 0.064 0.064 ;
END VIA78

VIA VIA67 Default
  LAYER M6 ;
    RECT -0.108 -0.064 0.108 0.064 ;
  LAYER M7 ;
    RECT -0.064 -0.108 0.064 0.108 ;
  LAYER V6 ;
    RECT -0.064 -0.064 0.064 0.064 ;
END VIA67

VIA VIA56 Default
  LAYER M5 ;
    RECT -0.048 -0.108 0.048 0.108 ;
  LAYER M6 ;
    RECT -0.092 -0.064 0.092 0.064 ;
  LAYER V5 ;
    RECT -0.048 -0.064 0.048 0.064 ;
END VIA56

VIA VIA45 Default
  LAYER M4 ;
    RECT -0.092 -0.048 0.092 0.048 ;
  LAYER M5 ;
    RECT -0.048 -0.092 0.048 0.092 ;
  LAYER V4 ;
    RECT -0.048 -0.048 0.048 0.048 ;
END VIA45

VIA VIA34 Default
  LAYER M3 ;
    RECT -0.036 -0.068 0.036 0.068 ;
  LAYER M4 ;
    RECT -0.080 -0.048 0.080 0.048 ;
  LAYER V3 ;
    RECT -0.036 -0.048 0.036 0.048 ;
END VIA34

VIA VIA23 Default
  LAYER M2 ;
    RECT -0.056 -0.036 0.056 0.036 ;
  LAYER M3 ;
    RECT -0.036 -0.056 0.036 0.056 ;
  LAYER V2 ;
    RECT -0.036 -0.036 0.036 0.036 ;
END VIA23

VIA VIA12 Default
  LAYER M1 ;
    RECT -0.036 -0.044 0.036 0.044 ;
  LAYER M2 ;
    RECT -0.056 -0.036 0.056 0.036 ;
  LAYER V1 ;
    RECT -0.036 -0.036 0.036 0.036 ;
END VIA12

#################################
### VIARULE GENERATE DEFAULTS ###
#################################

VIARULE Pad_M9 GENERATE DEFAULT
  LAYER M9 ;
    ENCLOSURE 0 0.0 ;
  LAYER Pad ;
    ENCLOSURE 0.044 0 ;
  LAYER V9 ;
    RECT -0.064 -0.064 0.064 0.064 ;
    SPACING 0.312 BY 0.312 ;
END Pad_M9

VIARULE M9_M8 GENERATE DEFAULT
  LAYER M8 ;
    ENCLOSURE 0.0 0 ;
  LAYER M9 ;
    ENCLOSURE 0 0.08 ;
  LAYER V8 ;
    RECT -0.08 -0.08 0.08 0.08 ;
    SPACING 0.388 BY 0.388 ;
END M9_M8

VIARULE M8_M7 GENERATE DEFAULT
  LAYER M7 ;
    ENCLOSURE 0.0 0.0 ;
  LAYER M8 ;
    ENCLOSURE 0.044 0 ;
  LAYER V7 ;
    RECT -0.064 -0.064 0.064 0.064 ;
    SPACING 0.312 BY 0.312 ;
END M8_M7

VIARULE M7_M6 GENERATE DEFAULT
  LAYER M6 ;
    ENCLOSURE 0.044 0 ;
  LAYER M7 ;
    ENCLOSURE 0 0.044 ;
  LAYER V6 ;
    RECT -0.064 -0.064 0.064 0.064 ;
    SPACING 0.312 BY 0.312 ;
END M7_M6

VIARULE M6_M5 GENERATE DEFAULT
  LAYER M5 ;
    ENCLOSURE 0.044 0.0 ;
    WIDTH 0.096 TO 0.096 ;
  LAYER M6 ;
    ENCLOSURE 0.044 0 ;
    WIDTH 0.128 TO 0.128 ;
  LAYER V5 ;
    RECT -0.048 -0.064 0.048 0.064 ;
    SPACING 0.232 BY 1.232 ;    # purposely crazy to avoid dual cut on routing
END M6_M5


# to make the wide vias for power stripes (still SAV)

VIARULE M3_M2widePWR0p936 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.0 0.0 ;
  LAYER M3 ;
    ENCLOSURE 0.0 0.0 ;
    WIDTH 0.936 TO 0.936 ;
  LAYER V2 ;
    RECT -0.468 -0.036 0.468 0.036 ;
    SPACING 1.108 BY 0.144 ;
END M3_M2widePWR0p936

# to make the wide vias for powers (still SAV)

VIARULE M4_M3widePWR0p864 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.0 0.0 ;
    WIDTH 0.934 TO 0.938 ;
  LAYER M4 ;
    ENCLOSURE 0.0 0.0 ;
    WIDTH 0.862 TO 0.866 ;
  LAYER V3 ;
    RECT -0.036 -0.432 0.036 0.432 ;
    SPACING 0.144 BY 1.108  ;
END M4_M3widePWR0p864

# to make the wide vias for powers (still SAV)

VIARULE M5_M4widePWR0p864 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.0 0.0 ;
  LAYER M5 ;
    ENCLOSURE 0.0 0.0 ;
    WIDTH 0.864 TO 0.864 ;
  LAYER V4 ;
    RECT -0.432 -0.048 0.432 0.048 ;
    SPACING 2.128 BY 0.384 ;
END M5_M4widePWR0p864

# to make the wide vias for powers (still SAV)

VIARULE M6_M5widePWR1p152 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.0 0.0 ;
  LAYER M6 ;
    ENCLOSURE 0.0 0.0 ;
    WIDTH 1.152 TO 1.152 ;
  LAYER V5 ;
    RECT -0.048 -0.576 0.048 0.576 ;
    SPACING 0.384 BY 1.528  ;
END M6_M5widePWR1p152

# to make the wide vias for powers (still SAV)

VIARULE M7_M6widePWR1p152 GENERATE
  LAYER M6 ;
    ENCLOSURE 0.0 0.0 ;
  LAYER M7 ;
    ENCLOSURE 0.0 0.0 ;
    WIDTH 1.152 TO 1.152 ;
  LAYER V6 ;
    RECT -0.576 -0.064 0.576 0.064 ;
    SPACING 2.128 BY 0.384 ;
END M7_M6widePWR1p152

VIARULE M2_M1 GENERATE DEFAULT
  LAYER M1 ;
    ENCLOSURE 0 0.0 ;		
  LAYER M2 ;
    ENCLOSURE 0.008 0.0 ;
  LAYER V1 ;
    RECT -0.036 -0.036 0.036 0.036 ;
    SPACING 0.144 BY 0.144 ;
END M2_M1

END LIBRARY
