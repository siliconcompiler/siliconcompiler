VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO heartbeat
  FOREIGN heartbeat ;


  SIZE 30.4 BY 30.4 ;
  CLASS BLOCK ;
  PIN clk
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.0
           10.115
           0.21000000000000002
           10.185 ;
    END
  END clk
  PIN nreset
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.0
           20.195
           0.21000000000000002
           20.265 ;
    END
  END nreset
  PIN out
    DIRECTION inout ;
    USE signal ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 30.189999999999998
           15.155
           30.4
           15.225 ;
    END
  END out


END heartbeat

END LIBRARY